`timescale 1ns / 1ps


module full_add(a,b,cin,cout,s);<br>
input a,b,cin;<br>
output s,cout;<br>
wire r,r1,r2;<br>
xor(s,a,b,cin);<br>
and(r,a,b);<br>
and(r1,b,cin);<br>
and(r2,a,cin);<br>
or(cout,r,r1,r2);<br>
endmodule<br>
module half_adder(input a,input b,output cout,output s);<br>
xor(s,a,b);<br>
and(cout,a,b);<br>
endmodule<br>
module jani(input [63:0]a,input [63:0]b,output [127:0]p);<br>

<br>
wire [63:0]andpr1;<br>
<br>
wire [63:0]andpr2;<br>
<br>
wire [63:0]andpr3;<br>
<br>
wire [63:0]andpr4;
<br><br>
wire [63:0]andpr5;
<br><br>
wire [63:0]andpr6;

wire [63:0]andpr7;

wire [63:0]andpr8;

wire [63:0]andpr9;

wire [63:0]andpr10;

wire [63:0]andpr11;

wire [63:0]andpr12;

wire [63:0]andpr13;

wire [63:0]andpr14;

wire [63:0]andpr15;

wire [63:0]andpr16;

wire [63:0]andpr17;

wire [63:0]andpr18;

wire [63:0]andpr19;

wire [63:0]andpr20;

wire [63:0]andpr21;

wire [63:0]andpr22;

wire [63:0]andpr23;

wire [63:0]andpr24;

wire [63:0]andpr25;

wire [63:0]andpr26;

wire [63:0]andpr27;

wire [63:0]andpr28;

wire [63:0]andpr29;

wire [63:0]andpr30;

wire [63:0]andpr31;

wire [63:0]andpr32;

wire [63:0]andpr33;

wire [63:0]andpr34;

wire [63:0]andpr35;

wire [63:0]andpr36;

wire [63:0]andpr37;

wire [63:0]andpr38;

wire [63:0]andpr39;

wire [63:0]andpr40;

wire [63:0]andpr41;

wire [63:0]andpr42;

wire [63:0]andpr43;

wire [63:0]andpr44;

wire [63:0]andpr45;

wire [63:0]andpr46;

wire [63:0]andpr47;

wire [63:0]andpr48;

wire [63:0]andpr49;

wire [63:0]andpr50;

wire [63:0]andpr51;

wire [63:0]andpr52;

wire [63:0]andpr53;

wire [63:0]andpr54;

wire [63:0]andpr55;

wire [63:0]andpr56;

wire [63:0]andpr57;

wire [63:0]andpr58;

wire [63:0]andpr59;

wire [63:0]andpr60;

wire [63:0]andpr61;

wire [63:0]andpr62;

wire [63:0]andpr63;

wire [63:0]andpr64;


wire [62:0]s1;
wire [63:0]c1;

wire [62:0]s2;
wire [63:0]c2;

wire [62:0]s3;
wire [63:0]c3;

wire [62:0]s4;
wire [63:0]c4;

wire [62:0]s5;
wire [63:0]c5;

wire [62:0]s6;
wire [63:0]c6;

wire [62:0]s7;
wire [63:0]c7;

wire [62:0]s8;
wire [63:0]c8;

wire [62:0]s9;
wire [63:0]c9;

wire [62:0]s10;
wire [63:0]c10;

wire [62:0]s11;
wire [63:0]c11;

wire [62:0]s12;
wire [63:0]c12;

wire [62:0]s13;
wire [63:0]c13;

wire [62:0]s14;
wire [63:0]c14;

wire [62:0]s15;
wire [63:0]c15;

wire [62:0]s16;
wire [63:0]c16;

wire [62:0]s17;
wire [63:0]c17;

wire [62:0]s18;
wire [63:0]c18;

wire [62:0]s19;
wire [63:0]c19;

wire [62:0]s20;
wire [63:0]c20;

wire [62:0]s21;
wire [63:0]c21;

wire [62:0]s22;
wire [63:0]c22;

wire [62:0]s23;
wire [63:0]c23;

wire [62:0]s24;
wire [63:0]c24;

wire [62:0]s25;
wire [63:0]c25;

wire [62:0]s26;
wire [63:0]c26;

wire [62:0]s27;
wire [63:0]c27;

wire [62:0]s28;
wire [63:0]c28;

wire [62:0]s29;
wire [63:0]c29;

wire [62:0]s30;
wire [63:0]c30;

wire [62:0]s31;
wire [63:0]c31;

wire [62:0]s32;
wire [63:0]c32;

wire [62:0]s33;
wire [63:0]c33;

wire [62:0]s34;
wire [63:0]c34;

wire [62:0]s35;
wire [63:0]c35;

wire [62:0]s36;
wire [63:0]c36;

wire [62:0]s37;
wire [63:0]c37;

wire [62:0]s38;
wire [63:0]c38;

wire [62:0]s39;
wire [63:0]c39;

wire [62:0]s40;
wire [63:0]c40;

wire [62:0]s41;
wire [63:0]c41;

wire [62:0]s42;
wire [63:0]c42;

wire [62:0]s43;
wire [63:0]c43;

wire [62:0]s44;
wire [63:0]c44;

wire [62:0]s45;
wire [63:0]c45;

wire [62:0]s46;
wire [63:0]c46;

wire [62:0]s47;
wire [63:0]c47;

wire [62:0]s48;
wire [63:0]c48;

wire [62:0]s49;
wire [63:0]c49;

wire [62:0]s50;
wire [63:0]c50;

wire [62:0]s51;
wire [63:0]c51;

wire [62:0]s52;
wire [63:0]c52;

wire [62:0]s53;
wire [63:0]c53;

wire [62:0]s54;
wire [63:0]c54;

wire [62:0]s55;
wire [63:0]c55;

wire [62:0]s56;
wire [63:0]c56;

wire [62:0]s57;
wire [63:0]c57;

wire [62:0]s58;
wire [63:0]c58;

wire [62:0]s59;
wire [63:0]c59;

wire [62:0]s60;
wire [63:0]c60;

wire [62:0]s61;
wire [63:0]c61;

wire [62:0]s62;
wire [63:0]c62;

wire [63:0]c63;
wire c;
wire [127:0]p;
wire [63:0]si;


    
        and(andpr1[0],b[0],a[0]);
        
    
        and(andpr1[1],b[0],a[1]);
        
    
        and(andpr1[2],b[0],a[2]);
        
    
        and(andpr1[3],b[0],a[3]);
        
    
        and(andpr1[4],b[0],a[4]);
        
    
        and(andpr1[5],b[0],a[5]);
        
    
        and(andpr1[6],b[0],a[6]);
        
    
        and(andpr1[7],b[0],a[7]);
        
    
        and(andpr1[8],b[0],a[8]);
        
    
        and(andpr1[9],b[0],a[9]);
        
    
        and(andpr1[10],b[0],a[10]);
        
    
        and(andpr1[11],b[0],a[11]);
        
    
        and(andpr1[12],b[0],a[12]);
        
    
        and(andpr1[13],b[0],a[13]);
        
    
        and(andpr1[14],b[0],a[14]);
        
    
        and(andpr1[15],b[0],a[15]);
        
    
        and(andpr1[16],b[0],a[16]);
        
    
        and(andpr1[17],b[0],a[17]);
        
    
        and(andpr1[18],b[0],a[18]);
        
    
        and(andpr1[19],b[0],a[19]);
        
    
        and(andpr1[20],b[0],a[20]);
        
    
        and(andpr1[21],b[0],a[21]);
        
    
        and(andpr1[22],b[0],a[22]);
        
    
        and(andpr1[23],b[0],a[23]);
        
    
        and(andpr1[24],b[0],a[24]);
        
    
        and(andpr1[25],b[0],a[25]);
        
    
        and(andpr1[26],b[0],a[26]);
        
    
        and(andpr1[27],b[0],a[27]);
        
    
        and(andpr1[28],b[0],a[28]);
        
    
        and(andpr1[29],b[0],a[29]);
        
    
        and(andpr1[30],b[0],a[30]);
        
    
        and(andpr1[31],b[0],a[31]);
        
    
        and(andpr1[32],b[0],a[32]);
        
    
        and(andpr1[33],b[0],a[33]);
        
    
        and(andpr1[34],b[0],a[34]);
        
    
        and(andpr1[35],b[0],a[35]);
        
    
        and(andpr1[36],b[0],a[36]);
        
    
        and(andpr1[37],b[0],a[37]);
        
    
        and(andpr1[38],b[0],a[38]);
        
    
        and(andpr1[39],b[0],a[39]);
        
    
        and(andpr1[40],b[0],a[40]);
        
    
        and(andpr1[41],b[0],a[41]);
        
    
        and(andpr1[42],b[0],a[42]);
        
    
        and(andpr1[43],b[0],a[43]);
        
    
        and(andpr1[44],b[0],a[44]);
        
    
        and(andpr1[45],b[0],a[45]);
        
    
        and(andpr1[46],b[0],a[46]);
        
    
        and(andpr1[47],b[0],a[47]);
        
    
        and(andpr1[48],b[0],a[48]);
        
    
        and(andpr1[49],b[0],a[49]);
        
    
        and(andpr1[50],b[0],a[50]);
        
    
        and(andpr1[51],b[0],a[51]);
        
    
        and(andpr1[52],b[0],a[52]);
        
    
        and(andpr1[53],b[0],a[53]);
        
    
        and(andpr1[54],b[0],a[54]);
        
    
        and(andpr1[55],b[0],a[55]);
        
    
        and(andpr1[56],b[0],a[56]);
        
    
        and(andpr1[57],b[0],a[57]);
        
    
        and(andpr1[58],b[0],a[58]);
        
    
        and(andpr1[59],b[0],a[59]);
        
    
        and(andpr1[60],b[0],a[60]);
        
    
        and(andpr1[61],b[0],a[61]);
        
    
        and(andpr1[62],b[0],a[62]);
        
    
        and(andpr1[63],b[0],a[63]);
        
    
    not(si[0],andpr1[63]);

    
        and(andpr2[0],b[1],a[0]);
        
    
        and(andpr2[1],b[1],a[1]);
        
    
        and(andpr2[2],b[1],a[2]);
        
    
        and(andpr2[3],b[1],a[3]);
        
    
        and(andpr2[4],b[1],a[4]);
        
    
        and(andpr2[5],b[1],a[5]);
        
    
        and(andpr2[6],b[1],a[6]);
        
    
        and(andpr2[7],b[1],a[7]);
        
    
        and(andpr2[8],b[1],a[8]);
        
    
        and(andpr2[9],b[1],a[9]);
        
    
        and(andpr2[10],b[1],a[10]);
        
    
        and(andpr2[11],b[1],a[11]);
        
    
        and(andpr2[12],b[1],a[12]);
        
    
        and(andpr2[13],b[1],a[13]);
        
    
        and(andpr2[14],b[1],a[14]);
        
    
        and(andpr2[15],b[1],a[15]);
        
    
        and(andpr2[16],b[1],a[16]);
        
    
        and(andpr2[17],b[1],a[17]);
        
    
        and(andpr2[18],b[1],a[18]);
        
    
        and(andpr2[19],b[1],a[19]);
        
    
        and(andpr2[20],b[1],a[20]);
        
    
        and(andpr2[21],b[1],a[21]);
        
    
        and(andpr2[22],b[1],a[22]);
        
    
        and(andpr2[23],b[1],a[23]);
        
    
        and(andpr2[24],b[1],a[24]);
        
    
        and(andpr2[25],b[1],a[25]);
        
    
        and(andpr2[26],b[1],a[26]);
        
    
        and(andpr2[27],b[1],a[27]);
        
    
        and(andpr2[28],b[1],a[28]);
        
    
        and(andpr2[29],b[1],a[29]);
        
    
        and(andpr2[30],b[1],a[30]);
        
    
        and(andpr2[31],b[1],a[31]);
        
    
        and(andpr2[32],b[1],a[32]);
        
    
        and(andpr2[33],b[1],a[33]);
        
    
        and(andpr2[34],b[1],a[34]);
        
    
        and(andpr2[35],b[1],a[35]);
        
    
        and(andpr2[36],b[1],a[36]);
        
    
        and(andpr2[37],b[1],a[37]);
        
    
        and(andpr2[38],b[1],a[38]);
        
    
        and(andpr2[39],b[1],a[39]);
        
    
        and(andpr2[40],b[1],a[40]);
        
    
        and(andpr2[41],b[1],a[41]);
        
    
        and(andpr2[42],b[1],a[42]);
        
    
        and(andpr2[43],b[1],a[43]);
        
    
        and(andpr2[44],b[1],a[44]);
        
    
        and(andpr2[45],b[1],a[45]);
        
    
        and(andpr2[46],b[1],a[46]);
        
    
        and(andpr2[47],b[1],a[47]);
        
    
        and(andpr2[48],b[1],a[48]);
        
    
        and(andpr2[49],b[1],a[49]);
        
    
        and(andpr2[50],b[1],a[50]);
        
    
        and(andpr2[51],b[1],a[51]);
        
    
        and(andpr2[52],b[1],a[52]);
        
    
        and(andpr2[53],b[1],a[53]);
        
    
        and(andpr2[54],b[1],a[54]);
        
    
        and(andpr2[55],b[1],a[55]);
        
    
        and(andpr2[56],b[1],a[56]);
        
    
        and(andpr2[57],b[1],a[57]);
        
    
        and(andpr2[58],b[1],a[58]);
        
    
        and(andpr2[59],b[1],a[59]);
        
    
        and(andpr2[60],b[1],a[60]);
        
    
        and(andpr2[61],b[1],a[61]);
        
    
        and(andpr2[62],b[1],a[62]);
        
    
        and(andpr2[63],b[1],a[63]);
        
    
    not(si[1],andpr2[63]);

    
        and(andpr3[0],b[2],a[0]);
        
    
        and(andpr3[1],b[2],a[1]);
        
    
        and(andpr3[2],b[2],a[2]);
        
    
        and(andpr3[3],b[2],a[3]);
        
    
        and(andpr3[4],b[2],a[4]);
        
    
        and(andpr3[5],b[2],a[5]);
        
    
        and(andpr3[6],b[2],a[6]);
        
    
        and(andpr3[7],b[2],a[7]);
        
    
        and(andpr3[8],b[2],a[8]);
        
    
        and(andpr3[9],b[2],a[9]);
        
    
        and(andpr3[10],b[2],a[10]);
        
    
        and(andpr3[11],b[2],a[11]);
        
    
        and(andpr3[12],b[2],a[12]);
        
    
        and(andpr3[13],b[2],a[13]);
        
    
        and(andpr3[14],b[2],a[14]);
        
    
        and(andpr3[15],b[2],a[15]);
        
    
        and(andpr3[16],b[2],a[16]);
        
    
        and(andpr3[17],b[2],a[17]);
        
    
        and(andpr3[18],b[2],a[18]);
        
    
        and(andpr3[19],b[2],a[19]);
        
    
        and(andpr3[20],b[2],a[20]);
        
    
        and(andpr3[21],b[2],a[21]);
        
    
        and(andpr3[22],b[2],a[22]);
        
    
        and(andpr3[23],b[2],a[23]);
        
    
        and(andpr3[24],b[2],a[24]);
        
    
        and(andpr3[25],b[2],a[25]);
        
    
        and(andpr3[26],b[2],a[26]);
        
    
        and(andpr3[27],b[2],a[27]);
        
    
        and(andpr3[28],b[2],a[28]);
        
    
        and(andpr3[29],b[2],a[29]);
        
    
        and(andpr3[30],b[2],a[30]);
        
    
        and(andpr3[31],b[2],a[31]);
        
    
        and(andpr3[32],b[2],a[32]);
        
    
        and(andpr3[33],b[2],a[33]);
        
    
        and(andpr3[34],b[2],a[34]);
        
    
        and(andpr3[35],b[2],a[35]);
        
    
        and(andpr3[36],b[2],a[36]);
        
    
        and(andpr3[37],b[2],a[37]);
        
    
        and(andpr3[38],b[2],a[38]);
        
    
        and(andpr3[39],b[2],a[39]);
        
    
        and(andpr3[40],b[2],a[40]);
        
    
        and(andpr3[41],b[2],a[41]);
        
    
        and(andpr3[42],b[2],a[42]);
        
    
        and(andpr3[43],b[2],a[43]);
        
    
        and(andpr3[44],b[2],a[44]);
        
    
        and(andpr3[45],b[2],a[45]);
        
    
        and(andpr3[46],b[2],a[46]);
        
    
        and(andpr3[47],b[2],a[47]);
        
    
        and(andpr3[48],b[2],a[48]);
        
    
        and(andpr3[49],b[2],a[49]);
        
    
        and(andpr3[50],b[2],a[50]);
        
    
        and(andpr3[51],b[2],a[51]);
        
    
        and(andpr3[52],b[2],a[52]);
        
    
        and(andpr3[53],b[2],a[53]);
        
    
        and(andpr3[54],b[2],a[54]);
        
    
        and(andpr3[55],b[2],a[55]);
        
    
        and(andpr3[56],b[2],a[56]);
        
    
        and(andpr3[57],b[2],a[57]);
        
    
        and(andpr3[58],b[2],a[58]);
        
    
        and(andpr3[59],b[2],a[59]);
        
    
        and(andpr3[60],b[2],a[60]);
        
    
        and(andpr3[61],b[2],a[61]);
        
    
        and(andpr3[62],b[2],a[62]);
        
    
        and(andpr3[63],b[2],a[63]);
        
    
    not(si[2],andpr3[63]);

    
        and(andpr4[0],b[3],a[0]);
        
    
        and(andpr4[1],b[3],a[1]);
        
    
        and(andpr4[2],b[3],a[2]);
        
    
        and(andpr4[3],b[3],a[3]);
        
    
        and(andpr4[4],b[3],a[4]);
        
    
        and(andpr4[5],b[3],a[5]);
        
    
        and(andpr4[6],b[3],a[6]);
        
    
        and(andpr4[7],b[3],a[7]);
        
    
        and(andpr4[8],b[3],a[8]);
        
    
        and(andpr4[9],b[3],a[9]);
        
    
        and(andpr4[10],b[3],a[10]);
        
    
        and(andpr4[11],b[3],a[11]);
        
    
        and(andpr4[12],b[3],a[12]);
        
    
        and(andpr4[13],b[3],a[13]);
        
    
        and(andpr4[14],b[3],a[14]);
        
    
        and(andpr4[15],b[3],a[15]);
        
    
        and(andpr4[16],b[3],a[16]);
        
    
        and(andpr4[17],b[3],a[17]);
        
    
        and(andpr4[18],b[3],a[18]);
        
    
        and(andpr4[19],b[3],a[19]);
        
    
        and(andpr4[20],b[3],a[20]);
        
    
        and(andpr4[21],b[3],a[21]);
        
    
        and(andpr4[22],b[3],a[22]);
        
    
        and(andpr4[23],b[3],a[23]);
        
    
        and(andpr4[24],b[3],a[24]);
        
    
        and(andpr4[25],b[3],a[25]);
        
    
        and(andpr4[26],b[3],a[26]);
        
    
        and(andpr4[27],b[3],a[27]);
        
    
        and(andpr4[28],b[3],a[28]);
        
    
        and(andpr4[29],b[3],a[29]);
        
    
        and(andpr4[30],b[3],a[30]);
        
    
        and(andpr4[31],b[3],a[31]);
        
    
        and(andpr4[32],b[3],a[32]);
        
    
        and(andpr4[33],b[3],a[33]);
        
    
        and(andpr4[34],b[3],a[34]);
        
    
        and(andpr4[35],b[3],a[35]);
        
    
        and(andpr4[36],b[3],a[36]);
        
    
        and(andpr4[37],b[3],a[37]);
        
    
        and(andpr4[38],b[3],a[38]);
        
    
        and(andpr4[39],b[3],a[39]);
        
    
        and(andpr4[40],b[3],a[40]);
        
    
        and(andpr4[41],b[3],a[41]);
        
    
        and(andpr4[42],b[3],a[42]);
        
    
        and(andpr4[43],b[3],a[43]);
        
    
        and(andpr4[44],b[3],a[44]);
        
    
        and(andpr4[45],b[3],a[45]);
        
    
        and(andpr4[46],b[3],a[46]);
        
    
        and(andpr4[47],b[3],a[47]);
        
    
        and(andpr4[48],b[3],a[48]);
        
    
        and(andpr4[49],b[3],a[49]);
        
    
        and(andpr4[50],b[3],a[50]);
        
    
        and(andpr4[51],b[3],a[51]);
        
    
        and(andpr4[52],b[3],a[52]);
        
    
        and(andpr4[53],b[3],a[53]);
        
    
        and(andpr4[54],b[3],a[54]);
        
    
        and(andpr4[55],b[3],a[55]);
        
    
        and(andpr4[56],b[3],a[56]);
        
    
        and(andpr4[57],b[3],a[57]);
        
    
        and(andpr4[58],b[3],a[58]);
        
    
        and(andpr4[59],b[3],a[59]);
        
    
        and(andpr4[60],b[3],a[60]);
        
    
        and(andpr4[61],b[3],a[61]);
        
    
        and(andpr4[62],b[3],a[62]);
        
    
        and(andpr4[63],b[3],a[63]);
        
    
    not(si[3],andpr4[63]);

    
        and(andpr5[0],b[4],a[0]);
        
    
        and(andpr5[1],b[4],a[1]);
        
    
        and(andpr5[2],b[4],a[2]);
        
    
        and(andpr5[3],b[4],a[3]);
        
    
        and(andpr5[4],b[4],a[4]);
        
    
        and(andpr5[5],b[4],a[5]);
        
    
        and(andpr5[6],b[4],a[6]);
        
    
        and(andpr5[7],b[4],a[7]);
        
    
        and(andpr5[8],b[4],a[8]);
        
    
        and(andpr5[9],b[4],a[9]);
        
    
        and(andpr5[10],b[4],a[10]);
        
    
        and(andpr5[11],b[4],a[11]);
        
    
        and(andpr5[12],b[4],a[12]);
        
    
        and(andpr5[13],b[4],a[13]);
        
    
        and(andpr5[14],b[4],a[14]);
        
    
        and(andpr5[15],b[4],a[15]);
        
    
        and(andpr5[16],b[4],a[16]);
        
    
        and(andpr5[17],b[4],a[17]);
        
    
        and(andpr5[18],b[4],a[18]);
        
    
        and(andpr5[19],b[4],a[19]);
        
    
        and(andpr5[20],b[4],a[20]);
        
    
        and(andpr5[21],b[4],a[21]);
        
    
        and(andpr5[22],b[4],a[22]);
        
    
        and(andpr5[23],b[4],a[23]);
        
    
        and(andpr5[24],b[4],a[24]);
        
    
        and(andpr5[25],b[4],a[25]);
        
    
        and(andpr5[26],b[4],a[26]);
        
    
        and(andpr5[27],b[4],a[27]);
        
    
        and(andpr5[28],b[4],a[28]);
        
    
        and(andpr5[29],b[4],a[29]);
        
    
        and(andpr5[30],b[4],a[30]);
        
    
        and(andpr5[31],b[4],a[31]);
        
    
        and(andpr5[32],b[4],a[32]);
        
    
        and(andpr5[33],b[4],a[33]);
        
    
        and(andpr5[34],b[4],a[34]);
        
    
        and(andpr5[35],b[4],a[35]);
        
    
        and(andpr5[36],b[4],a[36]);
        
    
        and(andpr5[37],b[4],a[37]);
        
    
        and(andpr5[38],b[4],a[38]);
        
    
        and(andpr5[39],b[4],a[39]);
        
    
        and(andpr5[40],b[4],a[40]);
        
    
        and(andpr5[41],b[4],a[41]);
        
    
        and(andpr5[42],b[4],a[42]);
        
    
        and(andpr5[43],b[4],a[43]);
        
    
        and(andpr5[44],b[4],a[44]);
        
    
        and(andpr5[45],b[4],a[45]);
        
    
        and(andpr5[46],b[4],a[46]);
        
    
        and(andpr5[47],b[4],a[47]);
        
    
        and(andpr5[48],b[4],a[48]);
        
    
        and(andpr5[49],b[4],a[49]);
        
    
        and(andpr5[50],b[4],a[50]);
        
    
        and(andpr5[51],b[4],a[51]);
        
    
        and(andpr5[52],b[4],a[52]);
        
    
        and(andpr5[53],b[4],a[53]);
        
    
        and(andpr5[54],b[4],a[54]);
        
    
        and(andpr5[55],b[4],a[55]);
        
    
        and(andpr5[56],b[4],a[56]);
        
    
        and(andpr5[57],b[4],a[57]);
        
    
        and(andpr5[58],b[4],a[58]);
        
    
        and(andpr5[59],b[4],a[59]);
        
    
        and(andpr5[60],b[4],a[60]);
        
    
        and(andpr5[61],b[4],a[61]);
        
    
        and(andpr5[62],b[4],a[62]);
        
    
        and(andpr5[63],b[4],a[63]);
        
    
    not(si[4],andpr5[63]);

    
        and(andpr6[0],b[5],a[0]);
        
    
        and(andpr6[1],b[5],a[1]);
        
    
        and(andpr6[2],b[5],a[2]);
        
    
        and(andpr6[3],b[5],a[3]);
        
    
        and(andpr6[4],b[5],a[4]);
        
    
        and(andpr6[5],b[5],a[5]);
        
    
        and(andpr6[6],b[5],a[6]);
        
    
        and(andpr6[7],b[5],a[7]);
        
    
        and(andpr6[8],b[5],a[8]);
        
    
        and(andpr6[9],b[5],a[9]);
        
    
        and(andpr6[10],b[5],a[10]);
        
    
        and(andpr6[11],b[5],a[11]);
        
    
        and(andpr6[12],b[5],a[12]);
        
    
        and(andpr6[13],b[5],a[13]);
        
    
        and(andpr6[14],b[5],a[14]);
        
    
        and(andpr6[15],b[5],a[15]);
        
    
        and(andpr6[16],b[5],a[16]);
        
    
        and(andpr6[17],b[5],a[17]);
        
    
        and(andpr6[18],b[5],a[18]);
        
    
        and(andpr6[19],b[5],a[19]);
        
    
        and(andpr6[20],b[5],a[20]);
        
    
        and(andpr6[21],b[5],a[21]);
        
    
        and(andpr6[22],b[5],a[22]);
        
    
        and(andpr6[23],b[5],a[23]);
        
    
        and(andpr6[24],b[5],a[24]);
        
    
        and(andpr6[25],b[5],a[25]);
        
    
        and(andpr6[26],b[5],a[26]);
        
    
        and(andpr6[27],b[5],a[27]);
        
    
        and(andpr6[28],b[5],a[28]);
        
    
        and(andpr6[29],b[5],a[29]);
        
    
        and(andpr6[30],b[5],a[30]);
        
    
        and(andpr6[31],b[5],a[31]);
        
    
        and(andpr6[32],b[5],a[32]);
        
    
        and(andpr6[33],b[5],a[33]);
        
    
        and(andpr6[34],b[5],a[34]);
        
    
        and(andpr6[35],b[5],a[35]);
        
    
        and(andpr6[36],b[5],a[36]);
        
    
        and(andpr6[37],b[5],a[37]);
        
    
        and(andpr6[38],b[5],a[38]);
        
    
        and(andpr6[39],b[5],a[39]);
        
    
        and(andpr6[40],b[5],a[40]);
        
    
        and(andpr6[41],b[5],a[41]);
        
    
        and(andpr6[42],b[5],a[42]);
        
    
        and(andpr6[43],b[5],a[43]);
        
    
        and(andpr6[44],b[5],a[44]);
        
    
        and(andpr6[45],b[5],a[45]);
        
    
        and(andpr6[46],b[5],a[46]);
        
    
        and(andpr6[47],b[5],a[47]);
        
    
        and(andpr6[48],b[5],a[48]);
        
    
        and(andpr6[49],b[5],a[49]);
        
    
        and(andpr6[50],b[5],a[50]);
        
    
        and(andpr6[51],b[5],a[51]);
        
    
        and(andpr6[52],b[5],a[52]);
        
    
        and(andpr6[53],b[5],a[53]);
        
    
        and(andpr6[54],b[5],a[54]);
        
    
        and(andpr6[55],b[5],a[55]);
        
    
        and(andpr6[56],b[5],a[56]);
        
    
        and(andpr6[57],b[5],a[57]);
        
    
        and(andpr6[58],b[5],a[58]);
        
    
        and(andpr6[59],b[5],a[59]);
        
    
        and(andpr6[60],b[5],a[60]);
        
    
        and(andpr6[61],b[5],a[61]);
        
    
        and(andpr6[62],b[5],a[62]);
        
    
        and(andpr6[63],b[5],a[63]);
        
    
    not(si[5],andpr6[63]);

    
        and(andpr7[0],b[6],a[0]);
        
    
        and(andpr7[1],b[6],a[1]);
        
    
        and(andpr7[2],b[6],a[2]);
        
    
        and(andpr7[3],b[6],a[3]);
        
    
        and(andpr7[4],b[6],a[4]);
        
    
        and(andpr7[5],b[6],a[5]);
        
    
        and(andpr7[6],b[6],a[6]);
        
    
        and(andpr7[7],b[6],a[7]);
        
    
        and(andpr7[8],b[6],a[8]);
        
    
        and(andpr7[9],b[6],a[9]);
        
    
        and(andpr7[10],b[6],a[10]);
        
    
        and(andpr7[11],b[6],a[11]);
        
    
        and(andpr7[12],b[6],a[12]);
        
    
        and(andpr7[13],b[6],a[13]);
        
    
        and(andpr7[14],b[6],a[14]);
        
    
        and(andpr7[15],b[6],a[15]);
        
    
        and(andpr7[16],b[6],a[16]);
        
    
        and(andpr7[17],b[6],a[17]);
        
    
        and(andpr7[18],b[6],a[18]);
        
    
        and(andpr7[19],b[6],a[19]);
        
    
        and(andpr7[20],b[6],a[20]);
        
    
        and(andpr7[21],b[6],a[21]);
        
    
        and(andpr7[22],b[6],a[22]);
        
    
        and(andpr7[23],b[6],a[23]);
        
    
        and(andpr7[24],b[6],a[24]);
        
    
        and(andpr7[25],b[6],a[25]);
        
    
        and(andpr7[26],b[6],a[26]);
        
    
        and(andpr7[27],b[6],a[27]);
        
    
        and(andpr7[28],b[6],a[28]);
        
    
        and(andpr7[29],b[6],a[29]);
        
    
        and(andpr7[30],b[6],a[30]);
        
    
        and(andpr7[31],b[6],a[31]);
        
    
        and(andpr7[32],b[6],a[32]);
        
    
        and(andpr7[33],b[6],a[33]);
        
    
        and(andpr7[34],b[6],a[34]);
        
    
        and(andpr7[35],b[6],a[35]);
        
    
        and(andpr7[36],b[6],a[36]);
        
    
        and(andpr7[37],b[6],a[37]);
        
    
        and(andpr7[38],b[6],a[38]);
        
    
        and(andpr7[39],b[6],a[39]);
        
    
        and(andpr7[40],b[6],a[40]);
        
    
        and(andpr7[41],b[6],a[41]);
        
    
        and(andpr7[42],b[6],a[42]);
        
    
        and(andpr7[43],b[6],a[43]);
        
    
        and(andpr7[44],b[6],a[44]);
        
    
        and(andpr7[45],b[6],a[45]);
        
    
        and(andpr7[46],b[6],a[46]);
        
    
        and(andpr7[47],b[6],a[47]);
        
    
        and(andpr7[48],b[6],a[48]);
        
    
        and(andpr7[49],b[6],a[49]);
        
    
        and(andpr7[50],b[6],a[50]);
        
    
        and(andpr7[51],b[6],a[51]);
        
    
        and(andpr7[52],b[6],a[52]);
        
    
        and(andpr7[53],b[6],a[53]);
        
    
        and(andpr7[54],b[6],a[54]);
        
    
        and(andpr7[55],b[6],a[55]);
        
    
        and(andpr7[56],b[6],a[56]);
        
    
        and(andpr7[57],b[6],a[57]);
        
    
        and(andpr7[58],b[6],a[58]);
        
    
        and(andpr7[59],b[6],a[59]);
        
    
        and(andpr7[60],b[6],a[60]);
        
    
        and(andpr7[61],b[6],a[61]);
        
    
        and(andpr7[62],b[6],a[62]);
        
    
        and(andpr7[63],b[6],a[63]);
        
    
    not(si[6],andpr7[63]);

    
        and(andpr8[0],b[7],a[0]);
        
    
        and(andpr8[1],b[7],a[1]);
        
    
        and(andpr8[2],b[7],a[2]);
        
    
        and(andpr8[3],b[7],a[3]);
        
    
        and(andpr8[4],b[7],a[4]);
        
    
        and(andpr8[5],b[7],a[5]);
        
    
        and(andpr8[6],b[7],a[6]);
        
    
        and(andpr8[7],b[7],a[7]);
        
    
        and(andpr8[8],b[7],a[8]);
        
    
        and(andpr8[9],b[7],a[9]);
        
    
        and(andpr8[10],b[7],a[10]);
        
    
        and(andpr8[11],b[7],a[11]);
        
    
        and(andpr8[12],b[7],a[12]);
        
    
        and(andpr8[13],b[7],a[13]);
        
    
        and(andpr8[14],b[7],a[14]);
        
    
        and(andpr8[15],b[7],a[15]);
        
    
        and(andpr8[16],b[7],a[16]);
        
    
        and(andpr8[17],b[7],a[17]);
        
    
        and(andpr8[18],b[7],a[18]);
        
    
        and(andpr8[19],b[7],a[19]);
        
    
        and(andpr8[20],b[7],a[20]);
        
    
        and(andpr8[21],b[7],a[21]);
        
    
        and(andpr8[22],b[7],a[22]);
        
    
        and(andpr8[23],b[7],a[23]);
        
    
        and(andpr8[24],b[7],a[24]);
        
    
        and(andpr8[25],b[7],a[25]);
        
    
        and(andpr8[26],b[7],a[26]);
        
    
        and(andpr8[27],b[7],a[27]);
        
    
        and(andpr8[28],b[7],a[28]);
        
    
        and(andpr8[29],b[7],a[29]);
        
    
        and(andpr8[30],b[7],a[30]);
        
    
        and(andpr8[31],b[7],a[31]);
        
    
        and(andpr8[32],b[7],a[32]);
        
    
        and(andpr8[33],b[7],a[33]);
        
    
        and(andpr8[34],b[7],a[34]);
        
    
        and(andpr8[35],b[7],a[35]);
        
    
        and(andpr8[36],b[7],a[36]);
        
    
        and(andpr8[37],b[7],a[37]);
        
    
        and(andpr8[38],b[7],a[38]);
        
    
        and(andpr8[39],b[7],a[39]);
        
    
        and(andpr8[40],b[7],a[40]);
        
    
        and(andpr8[41],b[7],a[41]);
        
    
        and(andpr8[42],b[7],a[42]);
        
    
        and(andpr8[43],b[7],a[43]);
        
    
        and(andpr8[44],b[7],a[44]);
        
    
        and(andpr8[45],b[7],a[45]);
        
    
        and(andpr8[46],b[7],a[46]);
        
    
        and(andpr8[47],b[7],a[47]);
        
    
        and(andpr8[48],b[7],a[48]);
        
    
        and(andpr8[49],b[7],a[49]);
        
    
        and(andpr8[50],b[7],a[50]);
        
    
        and(andpr8[51],b[7],a[51]);
        
    
        and(andpr8[52],b[7],a[52]);
        
    
        and(andpr8[53],b[7],a[53]);
        
    
        and(andpr8[54],b[7],a[54]);
        
    
        and(andpr8[55],b[7],a[55]);
        
    
        and(andpr8[56],b[7],a[56]);
        
    
        and(andpr8[57],b[7],a[57]);
        
    
        and(andpr8[58],b[7],a[58]);
        
    
        and(andpr8[59],b[7],a[59]);
        
    
        and(andpr8[60],b[7],a[60]);
        
    
        and(andpr8[61],b[7],a[61]);
        
    
        and(andpr8[62],b[7],a[62]);
        
    
        and(andpr8[63],b[7],a[63]);
        
    
    not(si[7],andpr8[63]);

    
        and(andpr9[0],b[8],a[0]);
        
    
        and(andpr9[1],b[8],a[1]);
        
    
        and(andpr9[2],b[8],a[2]);
        
    
        and(andpr9[3],b[8],a[3]);
        
    
        and(andpr9[4],b[8],a[4]);
        
    
        and(andpr9[5],b[8],a[5]);
        
    
        and(andpr9[6],b[8],a[6]);
        
    
        and(andpr9[7],b[8],a[7]);
        
    
        and(andpr9[8],b[8],a[8]);
        
    
        and(andpr9[9],b[8],a[9]);
        
    
        and(andpr9[10],b[8],a[10]);
        
    
        and(andpr9[11],b[8],a[11]);
        
    
        and(andpr9[12],b[8],a[12]);
        
    
        and(andpr9[13],b[8],a[13]);
        
    
        and(andpr9[14],b[8],a[14]);
        
    
        and(andpr9[15],b[8],a[15]);
        
    
        and(andpr9[16],b[8],a[16]);
        
    
        and(andpr9[17],b[8],a[17]);
        
    
        and(andpr9[18],b[8],a[18]);
        
    
        and(andpr9[19],b[8],a[19]);
        
    
        and(andpr9[20],b[8],a[20]);
        
    
        and(andpr9[21],b[8],a[21]);
        
    
        and(andpr9[22],b[8],a[22]);
        
    
        and(andpr9[23],b[8],a[23]);
        
    
        and(andpr9[24],b[8],a[24]);
        
    
        and(andpr9[25],b[8],a[25]);
        
    
        and(andpr9[26],b[8],a[26]);
        
    
        and(andpr9[27],b[8],a[27]);
        
    
        and(andpr9[28],b[8],a[28]);
        
    
        and(andpr9[29],b[8],a[29]);
        
    
        and(andpr9[30],b[8],a[30]);
        
    
        and(andpr9[31],b[8],a[31]);
        
    
        and(andpr9[32],b[8],a[32]);
        
    
        and(andpr9[33],b[8],a[33]);
        
    
        and(andpr9[34],b[8],a[34]);
        
    
        and(andpr9[35],b[8],a[35]);
        
    
        and(andpr9[36],b[8],a[36]);
        
    
        and(andpr9[37],b[8],a[37]);
        
    
        and(andpr9[38],b[8],a[38]);
        
    
        and(andpr9[39],b[8],a[39]);
        
    
        and(andpr9[40],b[8],a[40]);
        
    
        and(andpr9[41],b[8],a[41]);
        
    
        and(andpr9[42],b[8],a[42]);
        
    
        and(andpr9[43],b[8],a[43]);
        
    
        and(andpr9[44],b[8],a[44]);
        
    
        and(andpr9[45],b[8],a[45]);
        
    
        and(andpr9[46],b[8],a[46]);
        
    
        and(andpr9[47],b[8],a[47]);
        
    
        and(andpr9[48],b[8],a[48]);
        
    
        and(andpr9[49],b[8],a[49]);
        
    
        and(andpr9[50],b[8],a[50]);
        
    
        and(andpr9[51],b[8],a[51]);
        
    
        and(andpr9[52],b[8],a[52]);
        
    
        and(andpr9[53],b[8],a[53]);
        
    
        and(andpr9[54],b[8],a[54]);
        
    
        and(andpr9[55],b[8],a[55]);
        
    
        and(andpr9[56],b[8],a[56]);
        
    
        and(andpr9[57],b[8],a[57]);
        
    
        and(andpr9[58],b[8],a[58]);
        
    
        and(andpr9[59],b[8],a[59]);
        
    
        and(andpr9[60],b[8],a[60]);
        
    
        and(andpr9[61],b[8],a[61]);
        
    
        and(andpr9[62],b[8],a[62]);
        
    
        and(andpr9[63],b[8],a[63]);
        
    
    not(si[8],andpr9[63]);

    
        and(andpr10[0],b[9],a[0]);
        
    
        and(andpr10[1],b[9],a[1]);
        
    
        and(andpr10[2],b[9],a[2]);
        
    
        and(andpr10[3],b[9],a[3]);
        
    
        and(andpr10[4],b[9],a[4]);
        
    
        and(andpr10[5],b[9],a[5]);
        
    
        and(andpr10[6],b[9],a[6]);
        
    
        and(andpr10[7],b[9],a[7]);
        
    
        and(andpr10[8],b[9],a[8]);
        
    
        and(andpr10[9],b[9],a[9]);
        
    
        and(andpr10[10],b[9],a[10]);
        
    
        and(andpr10[11],b[9],a[11]);
        
    
        and(andpr10[12],b[9],a[12]);
        
    
        and(andpr10[13],b[9],a[13]);
        
    
        and(andpr10[14],b[9],a[14]);
        
    
        and(andpr10[15],b[9],a[15]);
        
    
        and(andpr10[16],b[9],a[16]);
        
    
        and(andpr10[17],b[9],a[17]);
        
    
        and(andpr10[18],b[9],a[18]);
        
    
        and(andpr10[19],b[9],a[19]);
        
    
        and(andpr10[20],b[9],a[20]);
        
    
        and(andpr10[21],b[9],a[21]);
        
    
        and(andpr10[22],b[9],a[22]);
        
    
        and(andpr10[23],b[9],a[23]);
        
    
        and(andpr10[24],b[9],a[24]);
        
    
        and(andpr10[25],b[9],a[25]);
        
    
        and(andpr10[26],b[9],a[26]);
        
    
        and(andpr10[27],b[9],a[27]);
        
    
        and(andpr10[28],b[9],a[28]);
        
    
        and(andpr10[29],b[9],a[29]);
        
    
        and(andpr10[30],b[9],a[30]);
        
    
        and(andpr10[31],b[9],a[31]);
        
    
        and(andpr10[32],b[9],a[32]);
        
    
        and(andpr10[33],b[9],a[33]);
        
    
        and(andpr10[34],b[9],a[34]);
        
    
        and(andpr10[35],b[9],a[35]);
        
    
        and(andpr10[36],b[9],a[36]);
        
    
        and(andpr10[37],b[9],a[37]);
        
    
        and(andpr10[38],b[9],a[38]);
        
    
        and(andpr10[39],b[9],a[39]);
        
    
        and(andpr10[40],b[9],a[40]);
        
    
        and(andpr10[41],b[9],a[41]);
        
    
        and(andpr10[42],b[9],a[42]);
        
    
        and(andpr10[43],b[9],a[43]);
        
    
        and(andpr10[44],b[9],a[44]);
        
    
        and(andpr10[45],b[9],a[45]);
        
    
        and(andpr10[46],b[9],a[46]);
        
    
        and(andpr10[47],b[9],a[47]);
        
    
        and(andpr10[48],b[9],a[48]);
        
    
        and(andpr10[49],b[9],a[49]);
        
    
        and(andpr10[50],b[9],a[50]);
        
    
        and(andpr10[51],b[9],a[51]);
        
    
        and(andpr10[52],b[9],a[52]);
        
    
        and(andpr10[53],b[9],a[53]);
        
    
        and(andpr10[54],b[9],a[54]);
        
    
        and(andpr10[55],b[9],a[55]);
        
    
        and(andpr10[56],b[9],a[56]);
        
    
        and(andpr10[57],b[9],a[57]);
        
    
        and(andpr10[58],b[9],a[58]);
        
    
        and(andpr10[59],b[9],a[59]);
        
    
        and(andpr10[60],b[9],a[60]);
        
    
        and(andpr10[61],b[9],a[61]);
        
    
        and(andpr10[62],b[9],a[62]);
        
    
        and(andpr10[63],b[9],a[63]);
        
    
    not(si[9],andpr10[63]);

    
        and(andpr11[0],b[10],a[0]);
        
    
        and(andpr11[1],b[10],a[1]);
        
    
        and(andpr11[2],b[10],a[2]);
        
    
        and(andpr11[3],b[10],a[3]);
        
    
        and(andpr11[4],b[10],a[4]);
        
    
        and(andpr11[5],b[10],a[5]);
        
    
        and(andpr11[6],b[10],a[6]);
        
    
        and(andpr11[7],b[10],a[7]);
        
    
        and(andpr11[8],b[10],a[8]);
        
    
        and(andpr11[9],b[10],a[9]);
        
    
        and(andpr11[10],b[10],a[10]);
        
    
        and(andpr11[11],b[10],a[11]);
        
    
        and(andpr11[12],b[10],a[12]);
        
    
        and(andpr11[13],b[10],a[13]);
        
    
        and(andpr11[14],b[10],a[14]);
        
    
        and(andpr11[15],b[10],a[15]);
        
    
        and(andpr11[16],b[10],a[16]);
        
    
        and(andpr11[17],b[10],a[17]);
        
    
        and(andpr11[18],b[10],a[18]);
        
    
        and(andpr11[19],b[10],a[19]);
        
    
        and(andpr11[20],b[10],a[20]);
        
    
        and(andpr11[21],b[10],a[21]);
        
    
        and(andpr11[22],b[10],a[22]);
        
    
        and(andpr11[23],b[10],a[23]);
        
    
        and(andpr11[24],b[10],a[24]);
        
    
        and(andpr11[25],b[10],a[25]);
        
    
        and(andpr11[26],b[10],a[26]);
        
    
        and(andpr11[27],b[10],a[27]);
        
    
        and(andpr11[28],b[10],a[28]);
        
    
        and(andpr11[29],b[10],a[29]);
        
    
        and(andpr11[30],b[10],a[30]);
        
    
        and(andpr11[31],b[10],a[31]);
        
    
        and(andpr11[32],b[10],a[32]);
        
    
        and(andpr11[33],b[10],a[33]);
        
    
        and(andpr11[34],b[10],a[34]);
        
    
        and(andpr11[35],b[10],a[35]);
        
    
        and(andpr11[36],b[10],a[36]);
        
    
        and(andpr11[37],b[10],a[37]);
        
    
        and(andpr11[38],b[10],a[38]);
        
    
        and(andpr11[39],b[10],a[39]);
        
    
        and(andpr11[40],b[10],a[40]);
        
    
        and(andpr11[41],b[10],a[41]);
        
    
        and(andpr11[42],b[10],a[42]);
        
    
        and(andpr11[43],b[10],a[43]);
        
    
        and(andpr11[44],b[10],a[44]);
        
    
        and(andpr11[45],b[10],a[45]);
        
    
        and(andpr11[46],b[10],a[46]);
        
    
        and(andpr11[47],b[10],a[47]);
        
    
        and(andpr11[48],b[10],a[48]);
        
    
        and(andpr11[49],b[10],a[49]);
        
    
        and(andpr11[50],b[10],a[50]);
        
    
        and(andpr11[51],b[10],a[51]);
        
    
        and(andpr11[52],b[10],a[52]);
        
    
        and(andpr11[53],b[10],a[53]);
        
    
        and(andpr11[54],b[10],a[54]);
        
    
        and(andpr11[55],b[10],a[55]);
        
    
        and(andpr11[56],b[10],a[56]);
        
    
        and(andpr11[57],b[10],a[57]);
        
    
        and(andpr11[58],b[10],a[58]);
        
    
        and(andpr11[59],b[10],a[59]);
        
    
        and(andpr11[60],b[10],a[60]);
        
    
        and(andpr11[61],b[10],a[61]);
        
    
        and(andpr11[62],b[10],a[62]);
        
    
        and(andpr11[63],b[10],a[63]);
        
    
    not(si[10],andpr11[63]);

    
        and(andpr12[0],b[11],a[0]);
        
    
        and(andpr12[1],b[11],a[1]);
        
    
        and(andpr12[2],b[11],a[2]);
        
    
        and(andpr12[3],b[11],a[3]);
        
    
        and(andpr12[4],b[11],a[4]);
        
    
        and(andpr12[5],b[11],a[5]);
        
    
        and(andpr12[6],b[11],a[6]);
        
    
        and(andpr12[7],b[11],a[7]);
        
    
        and(andpr12[8],b[11],a[8]);
        
    
        and(andpr12[9],b[11],a[9]);
        
    
        and(andpr12[10],b[11],a[10]);
        
    
        and(andpr12[11],b[11],a[11]);
        
    
        and(andpr12[12],b[11],a[12]);
        
    
        and(andpr12[13],b[11],a[13]);
        
    
        and(andpr12[14],b[11],a[14]);
        
    
        and(andpr12[15],b[11],a[15]);
        
    
        and(andpr12[16],b[11],a[16]);
        
    
        and(andpr12[17],b[11],a[17]);
        
    
        and(andpr12[18],b[11],a[18]);
        
    
        and(andpr12[19],b[11],a[19]);
        
    
        and(andpr12[20],b[11],a[20]);
        
    
        and(andpr12[21],b[11],a[21]);
        
    
        and(andpr12[22],b[11],a[22]);
        
    
        and(andpr12[23],b[11],a[23]);
        
    
        and(andpr12[24],b[11],a[24]);
        
    
        and(andpr12[25],b[11],a[25]);
        
    
        and(andpr12[26],b[11],a[26]);
        
    
        and(andpr12[27],b[11],a[27]);
        
    
        and(andpr12[28],b[11],a[28]);
        
    
        and(andpr12[29],b[11],a[29]);
        
    
        and(andpr12[30],b[11],a[30]);
        
    
        and(andpr12[31],b[11],a[31]);
        
    
        and(andpr12[32],b[11],a[32]);
        
    
        and(andpr12[33],b[11],a[33]);
        
    
        and(andpr12[34],b[11],a[34]);
        
    
        and(andpr12[35],b[11],a[35]);
        
    
        and(andpr12[36],b[11],a[36]);
        
    
        and(andpr12[37],b[11],a[37]);
        
    
        and(andpr12[38],b[11],a[38]);
        
    
        and(andpr12[39],b[11],a[39]);
        
    
        and(andpr12[40],b[11],a[40]);
        
    
        and(andpr12[41],b[11],a[41]);
        
    
        and(andpr12[42],b[11],a[42]);
        
    
        and(andpr12[43],b[11],a[43]);
        
    
        and(andpr12[44],b[11],a[44]);
        
    
        and(andpr12[45],b[11],a[45]);
        
    
        and(andpr12[46],b[11],a[46]);
        
    
        and(andpr12[47],b[11],a[47]);
        
    
        and(andpr12[48],b[11],a[48]);
        
    
        and(andpr12[49],b[11],a[49]);
        
    
        and(andpr12[50],b[11],a[50]);
        
    
        and(andpr12[51],b[11],a[51]);
        
    
        and(andpr12[52],b[11],a[52]);
        
    
        and(andpr12[53],b[11],a[53]);
        
    
        and(andpr12[54],b[11],a[54]);
        
    
        and(andpr12[55],b[11],a[55]);
        
    
        and(andpr12[56],b[11],a[56]);
        
    
        and(andpr12[57],b[11],a[57]);
        
    
        and(andpr12[58],b[11],a[58]);
        
    
        and(andpr12[59],b[11],a[59]);
        
    
        and(andpr12[60],b[11],a[60]);
        
    
        and(andpr12[61],b[11],a[61]);
        
    
        and(andpr12[62],b[11],a[62]);
        
    
        and(andpr12[63],b[11],a[63]);
        
    
    not(si[11],andpr12[63]);

    
        and(andpr13[0],b[12],a[0]);
        
    
        and(andpr13[1],b[12],a[1]);
        
    
        and(andpr13[2],b[12],a[2]);
        
    
        and(andpr13[3],b[12],a[3]);
        
    
        and(andpr13[4],b[12],a[4]);
        
    
        and(andpr13[5],b[12],a[5]);
        
    
        and(andpr13[6],b[12],a[6]);
        
    
        and(andpr13[7],b[12],a[7]);
        
    
        and(andpr13[8],b[12],a[8]);
        
    
        and(andpr13[9],b[12],a[9]);
        
    
        and(andpr13[10],b[12],a[10]);
        
    
        and(andpr13[11],b[12],a[11]);
        
    
        and(andpr13[12],b[12],a[12]);
        
    
        and(andpr13[13],b[12],a[13]);
        
    
        and(andpr13[14],b[12],a[14]);
        
    
        and(andpr13[15],b[12],a[15]);
        
    
        and(andpr13[16],b[12],a[16]);
        
    
        and(andpr13[17],b[12],a[17]);
        
    
        and(andpr13[18],b[12],a[18]);
        
    
        and(andpr13[19],b[12],a[19]);
        
    
        and(andpr13[20],b[12],a[20]);
        
    
        and(andpr13[21],b[12],a[21]);
        
    
        and(andpr13[22],b[12],a[22]);
        
    
        and(andpr13[23],b[12],a[23]);
        
    
        and(andpr13[24],b[12],a[24]);
        
    
        and(andpr13[25],b[12],a[25]);
        
    
        and(andpr13[26],b[12],a[26]);
        
    
        and(andpr13[27],b[12],a[27]);
        
    
        and(andpr13[28],b[12],a[28]);
        
    
        and(andpr13[29],b[12],a[29]);
        
    
        and(andpr13[30],b[12],a[30]);
        
    
        and(andpr13[31],b[12],a[31]);
        
    
        and(andpr13[32],b[12],a[32]);
        
    
        and(andpr13[33],b[12],a[33]);
        
    
        and(andpr13[34],b[12],a[34]);
        
    
        and(andpr13[35],b[12],a[35]);
        
    
        and(andpr13[36],b[12],a[36]);
        
    
        and(andpr13[37],b[12],a[37]);
        
    
        and(andpr13[38],b[12],a[38]);
        
    
        and(andpr13[39],b[12],a[39]);
        
    
        and(andpr13[40],b[12],a[40]);
        
    
        and(andpr13[41],b[12],a[41]);
        
    
        and(andpr13[42],b[12],a[42]);
        
    
        and(andpr13[43],b[12],a[43]);
        
    
        and(andpr13[44],b[12],a[44]);
        
    
        and(andpr13[45],b[12],a[45]);
        
    
        and(andpr13[46],b[12],a[46]);
        
    
        and(andpr13[47],b[12],a[47]);
        
    
        and(andpr13[48],b[12],a[48]);
        
    
        and(andpr13[49],b[12],a[49]);
        
    
        and(andpr13[50],b[12],a[50]);
        
    
        and(andpr13[51],b[12],a[51]);
        
    
        and(andpr13[52],b[12],a[52]);
        
    
        and(andpr13[53],b[12],a[53]);
        
    
        and(andpr13[54],b[12],a[54]);
        
    
        and(andpr13[55],b[12],a[55]);
        
    
        and(andpr13[56],b[12],a[56]);
        
    
        and(andpr13[57],b[12],a[57]);
        
    
        and(andpr13[58],b[12],a[58]);
        
    
        and(andpr13[59],b[12],a[59]);
        
    
        and(andpr13[60],b[12],a[60]);
        
    
        and(andpr13[61],b[12],a[61]);
        
    
        and(andpr13[62],b[12],a[62]);
        
    
        and(andpr13[63],b[12],a[63]);
        
    
    not(si[12],andpr13[63]);

    
        and(andpr14[0],b[13],a[0]);
        
    
        and(andpr14[1],b[13],a[1]);
        
    
        and(andpr14[2],b[13],a[2]);
        
    
        and(andpr14[3],b[13],a[3]);
        
    
        and(andpr14[4],b[13],a[4]);
        
    
        and(andpr14[5],b[13],a[5]);
        
    
        and(andpr14[6],b[13],a[6]);
        
    
        and(andpr14[7],b[13],a[7]);
        
    
        and(andpr14[8],b[13],a[8]);
        
    
        and(andpr14[9],b[13],a[9]);
        
    
        and(andpr14[10],b[13],a[10]);
        
    
        and(andpr14[11],b[13],a[11]);
        
    
        and(andpr14[12],b[13],a[12]);
        
    
        and(andpr14[13],b[13],a[13]);
        
    
        and(andpr14[14],b[13],a[14]);
        
    
        and(andpr14[15],b[13],a[15]);
        
    
        and(andpr14[16],b[13],a[16]);
        
    
        and(andpr14[17],b[13],a[17]);
        
    
        and(andpr14[18],b[13],a[18]);
        
    
        and(andpr14[19],b[13],a[19]);
        
    
        and(andpr14[20],b[13],a[20]);
        
    
        and(andpr14[21],b[13],a[21]);
        
    
        and(andpr14[22],b[13],a[22]);
        
    
        and(andpr14[23],b[13],a[23]);
        
    
        and(andpr14[24],b[13],a[24]);
        
    
        and(andpr14[25],b[13],a[25]);
        
    
        and(andpr14[26],b[13],a[26]);
        
    
        and(andpr14[27],b[13],a[27]);
        
    
        and(andpr14[28],b[13],a[28]);
        
    
        and(andpr14[29],b[13],a[29]);
        
    
        and(andpr14[30],b[13],a[30]);
        
    
        and(andpr14[31],b[13],a[31]);
        
    
        and(andpr14[32],b[13],a[32]);
        
    
        and(andpr14[33],b[13],a[33]);
        
    
        and(andpr14[34],b[13],a[34]);
        
    
        and(andpr14[35],b[13],a[35]);
        
    
        and(andpr14[36],b[13],a[36]);
        
    
        and(andpr14[37],b[13],a[37]);
        
    
        and(andpr14[38],b[13],a[38]);
        
    
        and(andpr14[39],b[13],a[39]);
        
    
        and(andpr14[40],b[13],a[40]);
        
    
        and(andpr14[41],b[13],a[41]);
        
    
        and(andpr14[42],b[13],a[42]);
        
    
        and(andpr14[43],b[13],a[43]);
        
    
        and(andpr14[44],b[13],a[44]);
        
    
        and(andpr14[45],b[13],a[45]);
        
    
        and(andpr14[46],b[13],a[46]);
        
    
        and(andpr14[47],b[13],a[47]);
        
    
        and(andpr14[48],b[13],a[48]);
        
    
        and(andpr14[49],b[13],a[49]);
        
    
        and(andpr14[50],b[13],a[50]);
        
    
        and(andpr14[51],b[13],a[51]);
        
    
        and(andpr14[52],b[13],a[52]);
        
    
        and(andpr14[53],b[13],a[53]);
        
    
        and(andpr14[54],b[13],a[54]);
        
    
        and(andpr14[55],b[13],a[55]);
        
    
        and(andpr14[56],b[13],a[56]);
        
    
        and(andpr14[57],b[13],a[57]);
        
    
        and(andpr14[58],b[13],a[58]);
        
    
        and(andpr14[59],b[13],a[59]);
        
    
        and(andpr14[60],b[13],a[60]);
        
    
        and(andpr14[61],b[13],a[61]);
        
    
        and(andpr14[62],b[13],a[62]);
        
    
        and(andpr14[63],b[13],a[63]);
        
    
    not(si[13],andpr14[63]);

    
        and(andpr15[0],b[14],a[0]);
        
    
        and(andpr15[1],b[14],a[1]);
        
    
        and(andpr15[2],b[14],a[2]);
        
    
        and(andpr15[3],b[14],a[3]);
        
    
        and(andpr15[4],b[14],a[4]);
        
    
        and(andpr15[5],b[14],a[5]);
        
    
        and(andpr15[6],b[14],a[6]);
        
    
        and(andpr15[7],b[14],a[7]);
        
    
        and(andpr15[8],b[14],a[8]);
        
    
        and(andpr15[9],b[14],a[9]);
        
    
        and(andpr15[10],b[14],a[10]);
        
    
        and(andpr15[11],b[14],a[11]);
        
    
        and(andpr15[12],b[14],a[12]);
        
    
        and(andpr15[13],b[14],a[13]);
        
    
        and(andpr15[14],b[14],a[14]);
        
    
        and(andpr15[15],b[14],a[15]);
        
    
        and(andpr15[16],b[14],a[16]);
        
    
        and(andpr15[17],b[14],a[17]);
        
    
        and(andpr15[18],b[14],a[18]);
        
    
        and(andpr15[19],b[14],a[19]);
        
    
        and(andpr15[20],b[14],a[20]);
        
    
        and(andpr15[21],b[14],a[21]);
        
    
        and(andpr15[22],b[14],a[22]);
        
    
        and(andpr15[23],b[14],a[23]);
        
    
        and(andpr15[24],b[14],a[24]);
        
    
        and(andpr15[25],b[14],a[25]);
        
    
        and(andpr15[26],b[14],a[26]);
        
    
        and(andpr15[27],b[14],a[27]);
        
    
        and(andpr15[28],b[14],a[28]);
        
    
        and(andpr15[29],b[14],a[29]);
        
    
        and(andpr15[30],b[14],a[30]);
        
    
        and(andpr15[31],b[14],a[31]);
        
    
        and(andpr15[32],b[14],a[32]);
        
    
        and(andpr15[33],b[14],a[33]);
        
    
        and(andpr15[34],b[14],a[34]);
        
    
        and(andpr15[35],b[14],a[35]);
        
    
        and(andpr15[36],b[14],a[36]);
        
    
        and(andpr15[37],b[14],a[37]);
        
    
        and(andpr15[38],b[14],a[38]);
        
    
        and(andpr15[39],b[14],a[39]);
        
    
        and(andpr15[40],b[14],a[40]);
        
    
        and(andpr15[41],b[14],a[41]);
        
    
        and(andpr15[42],b[14],a[42]);
        
    
        and(andpr15[43],b[14],a[43]);
        
    
        and(andpr15[44],b[14],a[44]);
        
    
        and(andpr15[45],b[14],a[45]);
        
    
        and(andpr15[46],b[14],a[46]);
        
    
        and(andpr15[47],b[14],a[47]);
        
    
        and(andpr15[48],b[14],a[48]);
        
    
        and(andpr15[49],b[14],a[49]);
        
    
        and(andpr15[50],b[14],a[50]);
        
    
        and(andpr15[51],b[14],a[51]);
        
    
        and(andpr15[52],b[14],a[52]);
        
    
        and(andpr15[53],b[14],a[53]);
        
    
        and(andpr15[54],b[14],a[54]);
        
    
        and(andpr15[55],b[14],a[55]);
        
    
        and(andpr15[56],b[14],a[56]);
        
    
        and(andpr15[57],b[14],a[57]);
        
    
        and(andpr15[58],b[14],a[58]);
        
    
        and(andpr15[59],b[14],a[59]);
        
    
        and(andpr15[60],b[14],a[60]);
        
    
        and(andpr15[61],b[14],a[61]);
        
    
        and(andpr15[62],b[14],a[62]);
        
    
        and(andpr15[63],b[14],a[63]);
        
    
    not(si[14],andpr15[63]);

    
        and(andpr16[0],b[15],a[0]);
        
    
        and(andpr16[1],b[15],a[1]);
        
    
        and(andpr16[2],b[15],a[2]);
        
    
        and(andpr16[3],b[15],a[3]);
        
    
        and(andpr16[4],b[15],a[4]);
        
    
        and(andpr16[5],b[15],a[5]);
        
    
        and(andpr16[6],b[15],a[6]);
        
    
        and(andpr16[7],b[15],a[7]);
        
    
        and(andpr16[8],b[15],a[8]);
        
    
        and(andpr16[9],b[15],a[9]);
        
    
        and(andpr16[10],b[15],a[10]);
        
    
        and(andpr16[11],b[15],a[11]);
        
    
        and(andpr16[12],b[15],a[12]);
        
    
        and(andpr16[13],b[15],a[13]);
        
    
        and(andpr16[14],b[15],a[14]);
        
    
        and(andpr16[15],b[15],a[15]);
        
    
        and(andpr16[16],b[15],a[16]);
        
    
        and(andpr16[17],b[15],a[17]);
        
    
        and(andpr16[18],b[15],a[18]);
        
    
        and(andpr16[19],b[15],a[19]);
        
    
        and(andpr16[20],b[15],a[20]);
        
    
        and(andpr16[21],b[15],a[21]);
        
    
        and(andpr16[22],b[15],a[22]);
        
    
        and(andpr16[23],b[15],a[23]);
        
    
        and(andpr16[24],b[15],a[24]);
        
    
        and(andpr16[25],b[15],a[25]);
        
    
        and(andpr16[26],b[15],a[26]);
        
    
        and(andpr16[27],b[15],a[27]);
        
    
        and(andpr16[28],b[15],a[28]);
        
    
        and(andpr16[29],b[15],a[29]);
        
    
        and(andpr16[30],b[15],a[30]);
        
    
        and(andpr16[31],b[15],a[31]);
        
    
        and(andpr16[32],b[15],a[32]);
        
    
        and(andpr16[33],b[15],a[33]);
        
    
        and(andpr16[34],b[15],a[34]);
        
    
        and(andpr16[35],b[15],a[35]);
        
    
        and(andpr16[36],b[15],a[36]);
        
    
        and(andpr16[37],b[15],a[37]);
        
    
        and(andpr16[38],b[15],a[38]);
        
    
        and(andpr16[39],b[15],a[39]);
        
    
        and(andpr16[40],b[15],a[40]);
        
    
        and(andpr16[41],b[15],a[41]);
        
    
        and(andpr16[42],b[15],a[42]);
        
    
        and(andpr16[43],b[15],a[43]);
        
    
        and(andpr16[44],b[15],a[44]);
        
    
        and(andpr16[45],b[15],a[45]);
        
    
        and(andpr16[46],b[15],a[46]);
        
    
        and(andpr16[47],b[15],a[47]);
        
    
        and(andpr16[48],b[15],a[48]);
        
    
        and(andpr16[49],b[15],a[49]);
        
    
        and(andpr16[50],b[15],a[50]);
        
    
        and(andpr16[51],b[15],a[51]);
        
    
        and(andpr16[52],b[15],a[52]);
        
    
        and(andpr16[53],b[15],a[53]);
        
    
        and(andpr16[54],b[15],a[54]);
        
    
        and(andpr16[55],b[15],a[55]);
        
    
        and(andpr16[56],b[15],a[56]);
        
    
        and(andpr16[57],b[15],a[57]);
        
    
        and(andpr16[58],b[15],a[58]);
        
    
        and(andpr16[59],b[15],a[59]);
        
    
        and(andpr16[60],b[15],a[60]);
        
    
        and(andpr16[61],b[15],a[61]);
        
    
        and(andpr16[62],b[15],a[62]);
        
    
        and(andpr16[63],b[15],a[63]);
        
    
    not(si[15],andpr16[63]);

    
        and(andpr17[0],b[16],a[0]);
        
    
        and(andpr17[1],b[16],a[1]);
        
    
        and(andpr17[2],b[16],a[2]);
        
    
        and(andpr17[3],b[16],a[3]);
        
    
        and(andpr17[4],b[16],a[4]);
        
    
        and(andpr17[5],b[16],a[5]);
        
    
        and(andpr17[6],b[16],a[6]);
        
    
        and(andpr17[7],b[16],a[7]);
        
    
        and(andpr17[8],b[16],a[8]);
        
    
        and(andpr17[9],b[16],a[9]);
        
    
        and(andpr17[10],b[16],a[10]);
        
    
        and(andpr17[11],b[16],a[11]);
        
    
        and(andpr17[12],b[16],a[12]);
        
    
        and(andpr17[13],b[16],a[13]);
        
    
        and(andpr17[14],b[16],a[14]);
        
    
        and(andpr17[15],b[16],a[15]);
        
    
        and(andpr17[16],b[16],a[16]);
        
    
        and(andpr17[17],b[16],a[17]);
        
    
        and(andpr17[18],b[16],a[18]);
        
    
        and(andpr17[19],b[16],a[19]);
        
    
        and(andpr17[20],b[16],a[20]);
        
    
        and(andpr17[21],b[16],a[21]);
        
    
        and(andpr17[22],b[16],a[22]);
        
    
        and(andpr17[23],b[16],a[23]);
        
    
        and(andpr17[24],b[16],a[24]);
        
    
        and(andpr17[25],b[16],a[25]);
        
    
        and(andpr17[26],b[16],a[26]);
        
    
        and(andpr17[27],b[16],a[27]);
        
    
        and(andpr17[28],b[16],a[28]);
        
    
        and(andpr17[29],b[16],a[29]);
        
    
        and(andpr17[30],b[16],a[30]);
        
    
        and(andpr17[31],b[16],a[31]);
        
    
        and(andpr17[32],b[16],a[32]);
        
    
        and(andpr17[33],b[16],a[33]);
        
    
        and(andpr17[34],b[16],a[34]);
        
    
        and(andpr17[35],b[16],a[35]);
        
    
        and(andpr17[36],b[16],a[36]);
        
    
        and(andpr17[37],b[16],a[37]);
        
    
        and(andpr17[38],b[16],a[38]);
        
    
        and(andpr17[39],b[16],a[39]);
        
    
        and(andpr17[40],b[16],a[40]);
        
    
        and(andpr17[41],b[16],a[41]);
        
    
        and(andpr17[42],b[16],a[42]);
        
    
        and(andpr17[43],b[16],a[43]);
        
    
        and(andpr17[44],b[16],a[44]);
        
    
        and(andpr17[45],b[16],a[45]);
        
    
        and(andpr17[46],b[16],a[46]);
        
    
        and(andpr17[47],b[16],a[47]);
        
    
        and(andpr17[48],b[16],a[48]);
        
    
        and(andpr17[49],b[16],a[49]);
        
    
        and(andpr17[50],b[16],a[50]);
        
    
        and(andpr17[51],b[16],a[51]);
        
    
        and(andpr17[52],b[16],a[52]);
        
    
        and(andpr17[53],b[16],a[53]);
        
    
        and(andpr17[54],b[16],a[54]);
        
    
        and(andpr17[55],b[16],a[55]);
        
    
        and(andpr17[56],b[16],a[56]);
        
    
        and(andpr17[57],b[16],a[57]);
        
    
        and(andpr17[58],b[16],a[58]);
        
    
        and(andpr17[59],b[16],a[59]);
        
    
        and(andpr17[60],b[16],a[60]);
        
    
        and(andpr17[61],b[16],a[61]);
        
    
        and(andpr17[62],b[16],a[62]);
        
    
        and(andpr17[63],b[16],a[63]);
        
    
    not(si[16],andpr17[63]);

    
        and(andpr18[0],b[17],a[0]);
        
    
        and(andpr18[1],b[17],a[1]);
        
    
        and(andpr18[2],b[17],a[2]);
        
    
        and(andpr18[3],b[17],a[3]);
        
    
        and(andpr18[4],b[17],a[4]);
        
    
        and(andpr18[5],b[17],a[5]);
        
    
        and(andpr18[6],b[17],a[6]);
        
    
        and(andpr18[7],b[17],a[7]);
        
    
        and(andpr18[8],b[17],a[8]);
        
    
        and(andpr18[9],b[17],a[9]);
        
    
        and(andpr18[10],b[17],a[10]);
        
    
        and(andpr18[11],b[17],a[11]);
        
    
        and(andpr18[12],b[17],a[12]);
        
    
        and(andpr18[13],b[17],a[13]);
        
    
        and(andpr18[14],b[17],a[14]);
        
    
        and(andpr18[15],b[17],a[15]);
        
    
        and(andpr18[16],b[17],a[16]);
        
    
        and(andpr18[17],b[17],a[17]);
        
    
        and(andpr18[18],b[17],a[18]);
        
    
        and(andpr18[19],b[17],a[19]);
        
    
        and(andpr18[20],b[17],a[20]);
        
    
        and(andpr18[21],b[17],a[21]);
        
    
        and(andpr18[22],b[17],a[22]);
        
    
        and(andpr18[23],b[17],a[23]);
        
    
        and(andpr18[24],b[17],a[24]);
        
    
        and(andpr18[25],b[17],a[25]);
        
    
        and(andpr18[26],b[17],a[26]);
        
    
        and(andpr18[27],b[17],a[27]);
        
    
        and(andpr18[28],b[17],a[28]);
        
    
        and(andpr18[29],b[17],a[29]);
        
    
        and(andpr18[30],b[17],a[30]);
        
    
        and(andpr18[31],b[17],a[31]);
        
    
        and(andpr18[32],b[17],a[32]);
        
    
        and(andpr18[33],b[17],a[33]);
        
    
        and(andpr18[34],b[17],a[34]);
        
    
        and(andpr18[35],b[17],a[35]);
        
    
        and(andpr18[36],b[17],a[36]);
        
    
        and(andpr18[37],b[17],a[37]);
        
    
        and(andpr18[38],b[17],a[38]);
        
    
        and(andpr18[39],b[17],a[39]);
        
    
        and(andpr18[40],b[17],a[40]);
        
    
        and(andpr18[41],b[17],a[41]);
        
    
        and(andpr18[42],b[17],a[42]);
        
    
        and(andpr18[43],b[17],a[43]);
        
    
        and(andpr18[44],b[17],a[44]);
        
    
        and(andpr18[45],b[17],a[45]);
        
    
        and(andpr18[46],b[17],a[46]);
        
    
        and(andpr18[47],b[17],a[47]);
        
    
        and(andpr18[48],b[17],a[48]);
        
    
        and(andpr18[49],b[17],a[49]);
        
    
        and(andpr18[50],b[17],a[50]);
        
    
        and(andpr18[51],b[17],a[51]);
        
    
        and(andpr18[52],b[17],a[52]);
        
    
        and(andpr18[53],b[17],a[53]);
        
    
        and(andpr18[54],b[17],a[54]);
        
    
        and(andpr18[55],b[17],a[55]);
        
    
        and(andpr18[56],b[17],a[56]);
        
    
        and(andpr18[57],b[17],a[57]);
        
    
        and(andpr18[58],b[17],a[58]);
        
    
        and(andpr18[59],b[17],a[59]);
        
    
        and(andpr18[60],b[17],a[60]);
        
    
        and(andpr18[61],b[17],a[61]);
        
    
        and(andpr18[62],b[17],a[62]);
        
    
        and(andpr18[63],b[17],a[63]);
        
    
    not(si[17],andpr18[63]);

    
        and(andpr19[0],b[18],a[0]);
        
    
        and(andpr19[1],b[18],a[1]);
        
    
        and(andpr19[2],b[18],a[2]);
        
    
        and(andpr19[3],b[18],a[3]);
        
    
        and(andpr19[4],b[18],a[4]);
        
    
        and(andpr19[5],b[18],a[5]);
        
    
        and(andpr19[6],b[18],a[6]);
        
    
        and(andpr19[7],b[18],a[7]);
        
    
        and(andpr19[8],b[18],a[8]);
        
    
        and(andpr19[9],b[18],a[9]);
        
    
        and(andpr19[10],b[18],a[10]);
        
    
        and(andpr19[11],b[18],a[11]);
        
    
        and(andpr19[12],b[18],a[12]);
        
    
        and(andpr19[13],b[18],a[13]);
        
    
        and(andpr19[14],b[18],a[14]);
        
    
        and(andpr19[15],b[18],a[15]);
        
    
        and(andpr19[16],b[18],a[16]);
        
    
        and(andpr19[17],b[18],a[17]);
        
    
        and(andpr19[18],b[18],a[18]);
        
    
        and(andpr19[19],b[18],a[19]);
        
    
        and(andpr19[20],b[18],a[20]);
        
    
        and(andpr19[21],b[18],a[21]);
        
    
        and(andpr19[22],b[18],a[22]);
        
    
        and(andpr19[23],b[18],a[23]);
        
    
        and(andpr19[24],b[18],a[24]);
        
    
        and(andpr19[25],b[18],a[25]);
        
    
        and(andpr19[26],b[18],a[26]);
        
    
        and(andpr19[27],b[18],a[27]);
        
    
        and(andpr19[28],b[18],a[28]);
        
    
        and(andpr19[29],b[18],a[29]);
        
    
        and(andpr19[30],b[18],a[30]);
        
    
        and(andpr19[31],b[18],a[31]);
        
    
        and(andpr19[32],b[18],a[32]);
        
    
        and(andpr19[33],b[18],a[33]);
        
    
        and(andpr19[34],b[18],a[34]);
        
    
        and(andpr19[35],b[18],a[35]);
        
    
        and(andpr19[36],b[18],a[36]);
        
    
        and(andpr19[37],b[18],a[37]);
        
    
        and(andpr19[38],b[18],a[38]);
        
    
        and(andpr19[39],b[18],a[39]);
        
    
        and(andpr19[40],b[18],a[40]);
        
    
        and(andpr19[41],b[18],a[41]);
        
    
        and(andpr19[42],b[18],a[42]);
        
    
        and(andpr19[43],b[18],a[43]);
        
    
        and(andpr19[44],b[18],a[44]);
        
    
        and(andpr19[45],b[18],a[45]);
        
    
        and(andpr19[46],b[18],a[46]);
        
    
        and(andpr19[47],b[18],a[47]);
        
    
        and(andpr19[48],b[18],a[48]);
        
    
        and(andpr19[49],b[18],a[49]);
        
    
        and(andpr19[50],b[18],a[50]);
        
    
        and(andpr19[51],b[18],a[51]);
        
    
        and(andpr19[52],b[18],a[52]);
        
    
        and(andpr19[53],b[18],a[53]);
        
    
        and(andpr19[54],b[18],a[54]);
        
    
        and(andpr19[55],b[18],a[55]);
        
    
        and(andpr19[56],b[18],a[56]);
        
    
        and(andpr19[57],b[18],a[57]);
        
    
        and(andpr19[58],b[18],a[58]);
        
    
        and(andpr19[59],b[18],a[59]);
        
    
        and(andpr19[60],b[18],a[60]);
        
    
        and(andpr19[61],b[18],a[61]);
        
    
        and(andpr19[62],b[18],a[62]);
        
    
        and(andpr19[63],b[18],a[63]);
        
    
    not(si[18],andpr19[63]);

    
        and(andpr20[0],b[19],a[0]);
        
    
        and(andpr20[1],b[19],a[1]);
        
    
        and(andpr20[2],b[19],a[2]);
        
    
        and(andpr20[3],b[19],a[3]);
        
    
        and(andpr20[4],b[19],a[4]);
        
    
        and(andpr20[5],b[19],a[5]);
        
    
        and(andpr20[6],b[19],a[6]);
        
    
        and(andpr20[7],b[19],a[7]);
        
    
        and(andpr20[8],b[19],a[8]);
        
    
        and(andpr20[9],b[19],a[9]);
        
    
        and(andpr20[10],b[19],a[10]);
        
    
        and(andpr20[11],b[19],a[11]);
        
    
        and(andpr20[12],b[19],a[12]);
        
    
        and(andpr20[13],b[19],a[13]);
        
    
        and(andpr20[14],b[19],a[14]);
        
    
        and(andpr20[15],b[19],a[15]);
        
    
        and(andpr20[16],b[19],a[16]);
        
    
        and(andpr20[17],b[19],a[17]);
        
    
        and(andpr20[18],b[19],a[18]);
        
    
        and(andpr20[19],b[19],a[19]);
        
    
        and(andpr20[20],b[19],a[20]);
        
    
        and(andpr20[21],b[19],a[21]);
        
    
        and(andpr20[22],b[19],a[22]);
        
    
        and(andpr20[23],b[19],a[23]);
        
    
        and(andpr20[24],b[19],a[24]);
        
    
        and(andpr20[25],b[19],a[25]);
        
    
        and(andpr20[26],b[19],a[26]);
        
    
        and(andpr20[27],b[19],a[27]);
        
    
        and(andpr20[28],b[19],a[28]);
        
    
        and(andpr20[29],b[19],a[29]);
        
    
        and(andpr20[30],b[19],a[30]);
        
    
        and(andpr20[31],b[19],a[31]);
        
    
        and(andpr20[32],b[19],a[32]);
        
    
        and(andpr20[33],b[19],a[33]);
        
    
        and(andpr20[34],b[19],a[34]);
        
    
        and(andpr20[35],b[19],a[35]);
        
    
        and(andpr20[36],b[19],a[36]);
        
    
        and(andpr20[37],b[19],a[37]);
        
    
        and(andpr20[38],b[19],a[38]);
        
    
        and(andpr20[39],b[19],a[39]);
        
    
        and(andpr20[40],b[19],a[40]);
        
    
        and(andpr20[41],b[19],a[41]);
        
    
        and(andpr20[42],b[19],a[42]);
        
    
        and(andpr20[43],b[19],a[43]);
        
    
        and(andpr20[44],b[19],a[44]);
        
    
        and(andpr20[45],b[19],a[45]);
        
    
        and(andpr20[46],b[19],a[46]);
        
    
        and(andpr20[47],b[19],a[47]);
        
    
        and(andpr20[48],b[19],a[48]);
        
    
        and(andpr20[49],b[19],a[49]);
        
    
        and(andpr20[50],b[19],a[50]);
        
    
        and(andpr20[51],b[19],a[51]);
        
    
        and(andpr20[52],b[19],a[52]);
        
    
        and(andpr20[53],b[19],a[53]);
        
    
        and(andpr20[54],b[19],a[54]);
        
    
        and(andpr20[55],b[19],a[55]);
        
    
        and(andpr20[56],b[19],a[56]);
        
    
        and(andpr20[57],b[19],a[57]);
        
    
        and(andpr20[58],b[19],a[58]);
        
    
        and(andpr20[59],b[19],a[59]);
        
    
        and(andpr20[60],b[19],a[60]);
        
    
        and(andpr20[61],b[19],a[61]);
        
    
        and(andpr20[62],b[19],a[62]);
        
    
        and(andpr20[63],b[19],a[63]);
        
    
    not(si[19],andpr20[63]);

    
        and(andpr21[0],b[20],a[0]);
        
    
        and(andpr21[1],b[20],a[1]);
        
    
        and(andpr21[2],b[20],a[2]);
        
    
        and(andpr21[3],b[20],a[3]);
        
    
        and(andpr21[4],b[20],a[4]);
        
    
        and(andpr21[5],b[20],a[5]);
        
    
        and(andpr21[6],b[20],a[6]);
        
    
        and(andpr21[7],b[20],a[7]);
        
    
        and(andpr21[8],b[20],a[8]);
        
    
        and(andpr21[9],b[20],a[9]);
        
    
        and(andpr21[10],b[20],a[10]);
        
    
        and(andpr21[11],b[20],a[11]);
        
    
        and(andpr21[12],b[20],a[12]);
        
    
        and(andpr21[13],b[20],a[13]);
        
    
        and(andpr21[14],b[20],a[14]);
        
    
        and(andpr21[15],b[20],a[15]);
        
    
        and(andpr21[16],b[20],a[16]);
        
    
        and(andpr21[17],b[20],a[17]);
        
    
        and(andpr21[18],b[20],a[18]);
        
    
        and(andpr21[19],b[20],a[19]);
        
    
        and(andpr21[20],b[20],a[20]);
        
    
        and(andpr21[21],b[20],a[21]);
        
    
        and(andpr21[22],b[20],a[22]);
        
    
        and(andpr21[23],b[20],a[23]);
        
    
        and(andpr21[24],b[20],a[24]);
        
    
        and(andpr21[25],b[20],a[25]);
        
    
        and(andpr21[26],b[20],a[26]);
        
    
        and(andpr21[27],b[20],a[27]);
        
    
        and(andpr21[28],b[20],a[28]);
        
    
        and(andpr21[29],b[20],a[29]);
        
    
        and(andpr21[30],b[20],a[30]);
        
    
        and(andpr21[31],b[20],a[31]);
        
    
        and(andpr21[32],b[20],a[32]);
        
    
        and(andpr21[33],b[20],a[33]);
        
    
        and(andpr21[34],b[20],a[34]);
        
    
        and(andpr21[35],b[20],a[35]);
        
    
        and(andpr21[36],b[20],a[36]);
        
    
        and(andpr21[37],b[20],a[37]);
        
    
        and(andpr21[38],b[20],a[38]);
        
    
        and(andpr21[39],b[20],a[39]);
        
    
        and(andpr21[40],b[20],a[40]);
        
    
        and(andpr21[41],b[20],a[41]);
        
    
        and(andpr21[42],b[20],a[42]);
        
    
        and(andpr21[43],b[20],a[43]);
        
    
        and(andpr21[44],b[20],a[44]);
        
    
        and(andpr21[45],b[20],a[45]);
        
    
        and(andpr21[46],b[20],a[46]);
        
    
        and(andpr21[47],b[20],a[47]);
        
    
        and(andpr21[48],b[20],a[48]);
        
    
        and(andpr21[49],b[20],a[49]);
        
    
        and(andpr21[50],b[20],a[50]);
        
    
        and(andpr21[51],b[20],a[51]);
        
    
        and(andpr21[52],b[20],a[52]);
        
    
        and(andpr21[53],b[20],a[53]);
        
    
        and(andpr21[54],b[20],a[54]);
        
    
        and(andpr21[55],b[20],a[55]);
        
    
        and(andpr21[56],b[20],a[56]);
        
    
        and(andpr21[57],b[20],a[57]);
        
    
        and(andpr21[58],b[20],a[58]);
        
    
        and(andpr21[59],b[20],a[59]);
        
    
        and(andpr21[60],b[20],a[60]);
        
    
        and(andpr21[61],b[20],a[61]);
        
    
        and(andpr21[62],b[20],a[62]);
        
    
        and(andpr21[63],b[20],a[63]);
        
    
    not(si[20],andpr21[63]);

    
        and(andpr22[0],b[21],a[0]);
        
    
        and(andpr22[1],b[21],a[1]);
        
    
        and(andpr22[2],b[21],a[2]);
        
    
        and(andpr22[3],b[21],a[3]);
        
    
        and(andpr22[4],b[21],a[4]);
        
    
        and(andpr22[5],b[21],a[5]);
        
    
        and(andpr22[6],b[21],a[6]);
        
    
        and(andpr22[7],b[21],a[7]);
        
    
        and(andpr22[8],b[21],a[8]);
        
    
        and(andpr22[9],b[21],a[9]);
        
    
        and(andpr22[10],b[21],a[10]);
        
    
        and(andpr22[11],b[21],a[11]);
        
    
        and(andpr22[12],b[21],a[12]);
        
    
        and(andpr22[13],b[21],a[13]);
        
    
        and(andpr22[14],b[21],a[14]);
        
    
        and(andpr22[15],b[21],a[15]);
        
    
        and(andpr22[16],b[21],a[16]);
        
    
        and(andpr22[17],b[21],a[17]);
        
    
        and(andpr22[18],b[21],a[18]);
        
    
        and(andpr22[19],b[21],a[19]);
        
    
        and(andpr22[20],b[21],a[20]);
        
    
        and(andpr22[21],b[21],a[21]);
        
    
        and(andpr22[22],b[21],a[22]);
        
    
        and(andpr22[23],b[21],a[23]);
        
    
        and(andpr22[24],b[21],a[24]);
        
    
        and(andpr22[25],b[21],a[25]);
        
    
        and(andpr22[26],b[21],a[26]);
        
    
        and(andpr22[27],b[21],a[27]);
        
    
        and(andpr22[28],b[21],a[28]);
        
    
        and(andpr22[29],b[21],a[29]);
        
    
        and(andpr22[30],b[21],a[30]);
        
    
        and(andpr22[31],b[21],a[31]);
        
    
        and(andpr22[32],b[21],a[32]);
        
    
        and(andpr22[33],b[21],a[33]);
        
    
        and(andpr22[34],b[21],a[34]);
        
    
        and(andpr22[35],b[21],a[35]);
        
    
        and(andpr22[36],b[21],a[36]);
        
    
        and(andpr22[37],b[21],a[37]);
        
    
        and(andpr22[38],b[21],a[38]);
        
    
        and(andpr22[39],b[21],a[39]);
        
    
        and(andpr22[40],b[21],a[40]);
        
    
        and(andpr22[41],b[21],a[41]);
        
    
        and(andpr22[42],b[21],a[42]);
        
    
        and(andpr22[43],b[21],a[43]);
        
    
        and(andpr22[44],b[21],a[44]);
        
    
        and(andpr22[45],b[21],a[45]);
        
    
        and(andpr22[46],b[21],a[46]);
        
    
        and(andpr22[47],b[21],a[47]);
        
    
        and(andpr22[48],b[21],a[48]);
        
    
        and(andpr22[49],b[21],a[49]);
        
    
        and(andpr22[50],b[21],a[50]);
        
    
        and(andpr22[51],b[21],a[51]);
        
    
        and(andpr22[52],b[21],a[52]);
        
    
        and(andpr22[53],b[21],a[53]);
        
    
        and(andpr22[54],b[21],a[54]);
        
    
        and(andpr22[55],b[21],a[55]);
        
    
        and(andpr22[56],b[21],a[56]);
        
    
        and(andpr22[57],b[21],a[57]);
        
    
        and(andpr22[58],b[21],a[58]);
        
    
        and(andpr22[59],b[21],a[59]);
        
    
        and(andpr22[60],b[21],a[60]);
        
    
        and(andpr22[61],b[21],a[61]);
        
    
        and(andpr22[62],b[21],a[62]);
        
    
        and(andpr22[63],b[21],a[63]);
        
    
    not(si[21],andpr22[63]);

    
        and(andpr23[0],b[22],a[0]);
        
    
        and(andpr23[1],b[22],a[1]);
        
    
        and(andpr23[2],b[22],a[2]);
        
    
        and(andpr23[3],b[22],a[3]);
        
    
        and(andpr23[4],b[22],a[4]);
        
    
        and(andpr23[5],b[22],a[5]);
        
    
        and(andpr23[6],b[22],a[6]);
        
    
        and(andpr23[7],b[22],a[7]);
        
    
        and(andpr23[8],b[22],a[8]);
        
    
        and(andpr23[9],b[22],a[9]);
        
    
        and(andpr23[10],b[22],a[10]);
        
    
        and(andpr23[11],b[22],a[11]);
        
    
        and(andpr23[12],b[22],a[12]);
        
    
        and(andpr23[13],b[22],a[13]);
        
    
        and(andpr23[14],b[22],a[14]);
        
    
        and(andpr23[15],b[22],a[15]);
        
    
        and(andpr23[16],b[22],a[16]);
        
    
        and(andpr23[17],b[22],a[17]);
        
    
        and(andpr23[18],b[22],a[18]);
        
    
        and(andpr23[19],b[22],a[19]);
        
    
        and(andpr23[20],b[22],a[20]);
        
    
        and(andpr23[21],b[22],a[21]);
        
    
        and(andpr23[22],b[22],a[22]);
        
    
        and(andpr23[23],b[22],a[23]);
        
    
        and(andpr23[24],b[22],a[24]);
        
    
        and(andpr23[25],b[22],a[25]);
        
    
        and(andpr23[26],b[22],a[26]);
        
    
        and(andpr23[27],b[22],a[27]);
        
    
        and(andpr23[28],b[22],a[28]);
        
    
        and(andpr23[29],b[22],a[29]);
        
    
        and(andpr23[30],b[22],a[30]);
        
    
        and(andpr23[31],b[22],a[31]);
        
    
        and(andpr23[32],b[22],a[32]);
        
    
        and(andpr23[33],b[22],a[33]);
        
    
        and(andpr23[34],b[22],a[34]);
        
    
        and(andpr23[35],b[22],a[35]);
        
    
        and(andpr23[36],b[22],a[36]);
        
    
        and(andpr23[37],b[22],a[37]);
        
    
        and(andpr23[38],b[22],a[38]);
        
    
        and(andpr23[39],b[22],a[39]);
        
    
        and(andpr23[40],b[22],a[40]);
        
    
        and(andpr23[41],b[22],a[41]);
        
    
        and(andpr23[42],b[22],a[42]);
        
    
        and(andpr23[43],b[22],a[43]);
        
    
        and(andpr23[44],b[22],a[44]);
        
    
        and(andpr23[45],b[22],a[45]);
        
    
        and(andpr23[46],b[22],a[46]);
        
    
        and(andpr23[47],b[22],a[47]);
        
    
        and(andpr23[48],b[22],a[48]);
        
    
        and(andpr23[49],b[22],a[49]);
        
    
        and(andpr23[50],b[22],a[50]);
        
    
        and(andpr23[51],b[22],a[51]);
        
    
        and(andpr23[52],b[22],a[52]);
        
    
        and(andpr23[53],b[22],a[53]);
        
    
        and(andpr23[54],b[22],a[54]);
        
    
        and(andpr23[55],b[22],a[55]);
        
    
        and(andpr23[56],b[22],a[56]);
        
    
        and(andpr23[57],b[22],a[57]);
        
    
        and(andpr23[58],b[22],a[58]);
        
    
        and(andpr23[59],b[22],a[59]);
        
    
        and(andpr23[60],b[22],a[60]);
        
    
        and(andpr23[61],b[22],a[61]);
        
    
        and(andpr23[62],b[22],a[62]);
        
    
        and(andpr23[63],b[22],a[63]);
        
    
    not(si[22],andpr23[63]);

    
        and(andpr24[0],b[23],a[0]);
        
    
        and(andpr24[1],b[23],a[1]);
        
    
        and(andpr24[2],b[23],a[2]);
        
    
        and(andpr24[3],b[23],a[3]);
        
    
        and(andpr24[4],b[23],a[4]);
        
    
        and(andpr24[5],b[23],a[5]);
        
    
        and(andpr24[6],b[23],a[6]);
        
    
        and(andpr24[7],b[23],a[7]);
        
    
        and(andpr24[8],b[23],a[8]);
        
    
        and(andpr24[9],b[23],a[9]);
        
    
        and(andpr24[10],b[23],a[10]);
        
    
        and(andpr24[11],b[23],a[11]);
        
    
        and(andpr24[12],b[23],a[12]);
        
    
        and(andpr24[13],b[23],a[13]);
        
    
        and(andpr24[14],b[23],a[14]);
        
    
        and(andpr24[15],b[23],a[15]);
        
    
        and(andpr24[16],b[23],a[16]);
        
    
        and(andpr24[17],b[23],a[17]);
        
    
        and(andpr24[18],b[23],a[18]);
        
    
        and(andpr24[19],b[23],a[19]);
        
    
        and(andpr24[20],b[23],a[20]);
        
    
        and(andpr24[21],b[23],a[21]);
        
    
        and(andpr24[22],b[23],a[22]);
        
    
        and(andpr24[23],b[23],a[23]);
        
    
        and(andpr24[24],b[23],a[24]);
        
    
        and(andpr24[25],b[23],a[25]);
        
    
        and(andpr24[26],b[23],a[26]);
        
    
        and(andpr24[27],b[23],a[27]);
        
    
        and(andpr24[28],b[23],a[28]);
        
    
        and(andpr24[29],b[23],a[29]);
        
    
        and(andpr24[30],b[23],a[30]);
        
    
        and(andpr24[31],b[23],a[31]);
        
    
        and(andpr24[32],b[23],a[32]);
        
    
        and(andpr24[33],b[23],a[33]);
        
    
        and(andpr24[34],b[23],a[34]);
        
    
        and(andpr24[35],b[23],a[35]);
        
    
        and(andpr24[36],b[23],a[36]);
        
    
        and(andpr24[37],b[23],a[37]);
        
    
        and(andpr24[38],b[23],a[38]);
        
    
        and(andpr24[39],b[23],a[39]);
        
    
        and(andpr24[40],b[23],a[40]);
        
    
        and(andpr24[41],b[23],a[41]);
        
    
        and(andpr24[42],b[23],a[42]);
        
    
        and(andpr24[43],b[23],a[43]);
        
    
        and(andpr24[44],b[23],a[44]);
        
    
        and(andpr24[45],b[23],a[45]);
        
    
        and(andpr24[46],b[23],a[46]);
        
    
        and(andpr24[47],b[23],a[47]);
        
    
        and(andpr24[48],b[23],a[48]);
        
    
        and(andpr24[49],b[23],a[49]);
        
    
        and(andpr24[50],b[23],a[50]);
        
    
        and(andpr24[51],b[23],a[51]);
        
    
        and(andpr24[52],b[23],a[52]);
        
    
        and(andpr24[53],b[23],a[53]);
        
    
        and(andpr24[54],b[23],a[54]);
        
    
        and(andpr24[55],b[23],a[55]);
        
    
        and(andpr24[56],b[23],a[56]);
        
    
        and(andpr24[57],b[23],a[57]);
        
    
        and(andpr24[58],b[23],a[58]);
        
    
        and(andpr24[59],b[23],a[59]);
        
    
        and(andpr24[60],b[23],a[60]);
        
    
        and(andpr24[61],b[23],a[61]);
        
    
        and(andpr24[62],b[23],a[62]);
        
    
        and(andpr24[63],b[23],a[63]);
        
    
    not(si[23],andpr24[63]);

    
        and(andpr25[0],b[24],a[0]);
        
    
        and(andpr25[1],b[24],a[1]);
        
    
        and(andpr25[2],b[24],a[2]);
        
    
        and(andpr25[3],b[24],a[3]);
        
    
        and(andpr25[4],b[24],a[4]);
        
    
        and(andpr25[5],b[24],a[5]);
        
    
        and(andpr25[6],b[24],a[6]);
        
    
        and(andpr25[7],b[24],a[7]);
        
    
        and(andpr25[8],b[24],a[8]);
        
    
        and(andpr25[9],b[24],a[9]);
        
    
        and(andpr25[10],b[24],a[10]);
        
    
        and(andpr25[11],b[24],a[11]);
        
    
        and(andpr25[12],b[24],a[12]);
        
    
        and(andpr25[13],b[24],a[13]);
        
    
        and(andpr25[14],b[24],a[14]);
        
    
        and(andpr25[15],b[24],a[15]);
        
    
        and(andpr25[16],b[24],a[16]);
        
    
        and(andpr25[17],b[24],a[17]);
        
    
        and(andpr25[18],b[24],a[18]);
        
    
        and(andpr25[19],b[24],a[19]);
        
    
        and(andpr25[20],b[24],a[20]);
        
    
        and(andpr25[21],b[24],a[21]);
        
    
        and(andpr25[22],b[24],a[22]);
        
    
        and(andpr25[23],b[24],a[23]);
        
    
        and(andpr25[24],b[24],a[24]);
        
    
        and(andpr25[25],b[24],a[25]);
        
    
        and(andpr25[26],b[24],a[26]);
        
    
        and(andpr25[27],b[24],a[27]);
        
    
        and(andpr25[28],b[24],a[28]);
        
    
        and(andpr25[29],b[24],a[29]);
        
    
        and(andpr25[30],b[24],a[30]);
        
    
        and(andpr25[31],b[24],a[31]);
        
    
        and(andpr25[32],b[24],a[32]);
        
    
        and(andpr25[33],b[24],a[33]);
        
    
        and(andpr25[34],b[24],a[34]);
        
    
        and(andpr25[35],b[24],a[35]);
        
    
        and(andpr25[36],b[24],a[36]);
        
    
        and(andpr25[37],b[24],a[37]);
        
    
        and(andpr25[38],b[24],a[38]);
        
    
        and(andpr25[39],b[24],a[39]);
        
    
        and(andpr25[40],b[24],a[40]);
        
    
        and(andpr25[41],b[24],a[41]);
        
    
        and(andpr25[42],b[24],a[42]);
        
    
        and(andpr25[43],b[24],a[43]);
        
    
        and(andpr25[44],b[24],a[44]);
        
    
        and(andpr25[45],b[24],a[45]);
        
    
        and(andpr25[46],b[24],a[46]);
        
    
        and(andpr25[47],b[24],a[47]);
        
    
        and(andpr25[48],b[24],a[48]);
        
    
        and(andpr25[49],b[24],a[49]);
        
    
        and(andpr25[50],b[24],a[50]);
        
    
        and(andpr25[51],b[24],a[51]);
        
    
        and(andpr25[52],b[24],a[52]);
        
    
        and(andpr25[53],b[24],a[53]);
        
    
        and(andpr25[54],b[24],a[54]);
        
    
        and(andpr25[55],b[24],a[55]);
        
    
        and(andpr25[56],b[24],a[56]);
        
    
        and(andpr25[57],b[24],a[57]);
        
    
        and(andpr25[58],b[24],a[58]);
        
    
        and(andpr25[59],b[24],a[59]);
        
    
        and(andpr25[60],b[24],a[60]);
        
    
        and(andpr25[61],b[24],a[61]);
        
    
        and(andpr25[62],b[24],a[62]);
        
    
        and(andpr25[63],b[24],a[63]);
        
    
    not(si[24],andpr25[63]);

    
        and(andpr26[0],b[25],a[0]);
        
    
        and(andpr26[1],b[25],a[1]);
        
    
        and(andpr26[2],b[25],a[2]);
        
    
        and(andpr26[3],b[25],a[3]);
        
    
        and(andpr26[4],b[25],a[4]);
        
    
        and(andpr26[5],b[25],a[5]);
        
    
        and(andpr26[6],b[25],a[6]);
        
    
        and(andpr26[7],b[25],a[7]);
        
    
        and(andpr26[8],b[25],a[8]);
        
    
        and(andpr26[9],b[25],a[9]);
        
    
        and(andpr26[10],b[25],a[10]);
        
    
        and(andpr26[11],b[25],a[11]);
        
    
        and(andpr26[12],b[25],a[12]);
        
    
        and(andpr26[13],b[25],a[13]);
        
    
        and(andpr26[14],b[25],a[14]);
        
    
        and(andpr26[15],b[25],a[15]);
        
    
        and(andpr26[16],b[25],a[16]);
        
    
        and(andpr26[17],b[25],a[17]);
        
    
        and(andpr26[18],b[25],a[18]);
        
    
        and(andpr26[19],b[25],a[19]);
        
    
        and(andpr26[20],b[25],a[20]);
        
    
        and(andpr26[21],b[25],a[21]);
        
    
        and(andpr26[22],b[25],a[22]);
        
    
        and(andpr26[23],b[25],a[23]);
        
    
        and(andpr26[24],b[25],a[24]);
        
    
        and(andpr26[25],b[25],a[25]);
        
    
        and(andpr26[26],b[25],a[26]);
        
    
        and(andpr26[27],b[25],a[27]);
        
    
        and(andpr26[28],b[25],a[28]);
        
    
        and(andpr26[29],b[25],a[29]);
        
    
        and(andpr26[30],b[25],a[30]);
        
    
        and(andpr26[31],b[25],a[31]);
        
    
        and(andpr26[32],b[25],a[32]);
        
    
        and(andpr26[33],b[25],a[33]);
        
    
        and(andpr26[34],b[25],a[34]);
        
    
        and(andpr26[35],b[25],a[35]);
        
    
        and(andpr26[36],b[25],a[36]);
        
    
        and(andpr26[37],b[25],a[37]);
        
    
        and(andpr26[38],b[25],a[38]);
        
    
        and(andpr26[39],b[25],a[39]);
        
    
        and(andpr26[40],b[25],a[40]);
        
    
        and(andpr26[41],b[25],a[41]);
        
    
        and(andpr26[42],b[25],a[42]);
        
    
        and(andpr26[43],b[25],a[43]);
        
    
        and(andpr26[44],b[25],a[44]);
        
    
        and(andpr26[45],b[25],a[45]);
        
    
        and(andpr26[46],b[25],a[46]);
        
    
        and(andpr26[47],b[25],a[47]);
        
    
        and(andpr26[48],b[25],a[48]);
        
    
        and(andpr26[49],b[25],a[49]);
        
    
        and(andpr26[50],b[25],a[50]);
        
    
        and(andpr26[51],b[25],a[51]);
        
    
        and(andpr26[52],b[25],a[52]);
        
    
        and(andpr26[53],b[25],a[53]);
        
    
        and(andpr26[54],b[25],a[54]);
        
    
        and(andpr26[55],b[25],a[55]);
        
    
        and(andpr26[56],b[25],a[56]);
        
    
        and(andpr26[57],b[25],a[57]);
        
    
        and(andpr26[58],b[25],a[58]);
        
    
        and(andpr26[59],b[25],a[59]);
        
    
        and(andpr26[60],b[25],a[60]);
        
    
        and(andpr26[61],b[25],a[61]);
        
    
        and(andpr26[62],b[25],a[62]);
        
    
        and(andpr26[63],b[25],a[63]);
        
    
    not(si[25],andpr26[63]);

    
        and(andpr27[0],b[26],a[0]);
        
    
        and(andpr27[1],b[26],a[1]);
        
    
        and(andpr27[2],b[26],a[2]);
        
    
        and(andpr27[3],b[26],a[3]);
        
    
        and(andpr27[4],b[26],a[4]);
        
    
        and(andpr27[5],b[26],a[5]);
        
    
        and(andpr27[6],b[26],a[6]);
        
    
        and(andpr27[7],b[26],a[7]);
        
    
        and(andpr27[8],b[26],a[8]);
        
    
        and(andpr27[9],b[26],a[9]);
        
    
        and(andpr27[10],b[26],a[10]);
        
    
        and(andpr27[11],b[26],a[11]);
        
    
        and(andpr27[12],b[26],a[12]);
        
    
        and(andpr27[13],b[26],a[13]);
        
    
        and(andpr27[14],b[26],a[14]);
        
    
        and(andpr27[15],b[26],a[15]);
        
    
        and(andpr27[16],b[26],a[16]);
        
    
        and(andpr27[17],b[26],a[17]);
        
    
        and(andpr27[18],b[26],a[18]);
        
    
        and(andpr27[19],b[26],a[19]);
        
    
        and(andpr27[20],b[26],a[20]);
        
    
        and(andpr27[21],b[26],a[21]);
        
    
        and(andpr27[22],b[26],a[22]);
        
    
        and(andpr27[23],b[26],a[23]);
        
    
        and(andpr27[24],b[26],a[24]);
        
    
        and(andpr27[25],b[26],a[25]);
        
    
        and(andpr27[26],b[26],a[26]);
        
    
        and(andpr27[27],b[26],a[27]);
        
    
        and(andpr27[28],b[26],a[28]);
        
    
        and(andpr27[29],b[26],a[29]);
        
    
        and(andpr27[30],b[26],a[30]);
        
    
        and(andpr27[31],b[26],a[31]);
        
    
        and(andpr27[32],b[26],a[32]);
        
    
        and(andpr27[33],b[26],a[33]);
        
    
        and(andpr27[34],b[26],a[34]);
        
    
        and(andpr27[35],b[26],a[35]);
        
    
        and(andpr27[36],b[26],a[36]);
        
    
        and(andpr27[37],b[26],a[37]);
        
    
        and(andpr27[38],b[26],a[38]);
        
    
        and(andpr27[39],b[26],a[39]);
        
    
        and(andpr27[40],b[26],a[40]);
        
    
        and(andpr27[41],b[26],a[41]);
        
    
        and(andpr27[42],b[26],a[42]);
        
    
        and(andpr27[43],b[26],a[43]);
        
    
        and(andpr27[44],b[26],a[44]);
        
    
        and(andpr27[45],b[26],a[45]);
        
    
        and(andpr27[46],b[26],a[46]);
        
    
        and(andpr27[47],b[26],a[47]);
        
    
        and(andpr27[48],b[26],a[48]);
        
    
        and(andpr27[49],b[26],a[49]);
        
    
        and(andpr27[50],b[26],a[50]);
        
    
        and(andpr27[51],b[26],a[51]);
        
    
        and(andpr27[52],b[26],a[52]);
        
    
        and(andpr27[53],b[26],a[53]);
        
    
        and(andpr27[54],b[26],a[54]);
        
    
        and(andpr27[55],b[26],a[55]);
        
    
        and(andpr27[56],b[26],a[56]);
        
    
        and(andpr27[57],b[26],a[57]);
        
    
        and(andpr27[58],b[26],a[58]);
        
    
        and(andpr27[59],b[26],a[59]);
        
    
        and(andpr27[60],b[26],a[60]);
        
    
        and(andpr27[61],b[26],a[61]);
        
    
        and(andpr27[62],b[26],a[62]);
        
    
        and(andpr27[63],b[26],a[63]);
        
    
    not(si[26],andpr27[63]);

    
        and(andpr28[0],b[27],a[0]);
        
    
        and(andpr28[1],b[27],a[1]);
        
    
        and(andpr28[2],b[27],a[2]);
        
    
        and(andpr28[3],b[27],a[3]);
        
    
        and(andpr28[4],b[27],a[4]);
        
    
        and(andpr28[5],b[27],a[5]);
        
    
        and(andpr28[6],b[27],a[6]);
        
    
        and(andpr28[7],b[27],a[7]);
        
    
        and(andpr28[8],b[27],a[8]);
        
    
        and(andpr28[9],b[27],a[9]);
        
    
        and(andpr28[10],b[27],a[10]);
        
    
        and(andpr28[11],b[27],a[11]);
        
    
        and(andpr28[12],b[27],a[12]);
        
    
        and(andpr28[13],b[27],a[13]);
        
    
        and(andpr28[14],b[27],a[14]);
        
    
        and(andpr28[15],b[27],a[15]);
        
    
        and(andpr28[16],b[27],a[16]);
        
    
        and(andpr28[17],b[27],a[17]);
        
    
        and(andpr28[18],b[27],a[18]);
        
    
        and(andpr28[19],b[27],a[19]);
        
    
        and(andpr28[20],b[27],a[20]);
        
    
        and(andpr28[21],b[27],a[21]);
        
    
        and(andpr28[22],b[27],a[22]);
        
    
        and(andpr28[23],b[27],a[23]);
        
    
        and(andpr28[24],b[27],a[24]);
        
    
        and(andpr28[25],b[27],a[25]);
        
    
        and(andpr28[26],b[27],a[26]);
        
    
        and(andpr28[27],b[27],a[27]);
        
    
        and(andpr28[28],b[27],a[28]);
        
    
        and(andpr28[29],b[27],a[29]);
        
    
        and(andpr28[30],b[27],a[30]);
        
    
        and(andpr28[31],b[27],a[31]);
        
    
        and(andpr28[32],b[27],a[32]);
        
    
        and(andpr28[33],b[27],a[33]);
        
    
        and(andpr28[34],b[27],a[34]);
        
    
        and(andpr28[35],b[27],a[35]);
        
    
        and(andpr28[36],b[27],a[36]);
        
    
        and(andpr28[37],b[27],a[37]);
        
    
        and(andpr28[38],b[27],a[38]);
        
    
        and(andpr28[39],b[27],a[39]);
        
    
        and(andpr28[40],b[27],a[40]);
        
    
        and(andpr28[41],b[27],a[41]);
        
    
        and(andpr28[42],b[27],a[42]);
        
    
        and(andpr28[43],b[27],a[43]);
        
    
        and(andpr28[44],b[27],a[44]);
        
    
        and(andpr28[45],b[27],a[45]);
        
    
        and(andpr28[46],b[27],a[46]);
        
    
        and(andpr28[47],b[27],a[47]);
        
    
        and(andpr28[48],b[27],a[48]);
        
    
        and(andpr28[49],b[27],a[49]);
        
    
        and(andpr28[50],b[27],a[50]);
        
    
        and(andpr28[51],b[27],a[51]);
        
    
        and(andpr28[52],b[27],a[52]);
        
    
        and(andpr28[53],b[27],a[53]);
        
    
        and(andpr28[54],b[27],a[54]);
        
    
        and(andpr28[55],b[27],a[55]);
        
    
        and(andpr28[56],b[27],a[56]);
        
    
        and(andpr28[57],b[27],a[57]);
        
    
        and(andpr28[58],b[27],a[58]);
        
    
        and(andpr28[59],b[27],a[59]);
        
    
        and(andpr28[60],b[27],a[60]);
        
    
        and(andpr28[61],b[27],a[61]);
        
    
        and(andpr28[62],b[27],a[62]);
        
    
        and(andpr28[63],b[27],a[63]);
        
    
    not(si[27],andpr28[63]);

    
        and(andpr29[0],b[28],a[0]);
        
    
        and(andpr29[1],b[28],a[1]);
        
    
        and(andpr29[2],b[28],a[2]);
        
    
        and(andpr29[3],b[28],a[3]);
        
    
        and(andpr29[4],b[28],a[4]);
        
    
        and(andpr29[5],b[28],a[5]);
        
    
        and(andpr29[6],b[28],a[6]);
        
    
        and(andpr29[7],b[28],a[7]);
        
    
        and(andpr29[8],b[28],a[8]);
        
    
        and(andpr29[9],b[28],a[9]);
        
    
        and(andpr29[10],b[28],a[10]);
        
    
        and(andpr29[11],b[28],a[11]);
        
    
        and(andpr29[12],b[28],a[12]);
        
    
        and(andpr29[13],b[28],a[13]);
        
    
        and(andpr29[14],b[28],a[14]);
        
    
        and(andpr29[15],b[28],a[15]);
        
    
        and(andpr29[16],b[28],a[16]);
        
    
        and(andpr29[17],b[28],a[17]);
        
    
        and(andpr29[18],b[28],a[18]);
        
    
        and(andpr29[19],b[28],a[19]);
        
    
        and(andpr29[20],b[28],a[20]);
        
    
        and(andpr29[21],b[28],a[21]);
        
    
        and(andpr29[22],b[28],a[22]);
        
    
        and(andpr29[23],b[28],a[23]);
        
    
        and(andpr29[24],b[28],a[24]);
        
    
        and(andpr29[25],b[28],a[25]);
        
    
        and(andpr29[26],b[28],a[26]);
        
    
        and(andpr29[27],b[28],a[27]);
        
    
        and(andpr29[28],b[28],a[28]);
        
    
        and(andpr29[29],b[28],a[29]);
        
    
        and(andpr29[30],b[28],a[30]);
        
    
        and(andpr29[31],b[28],a[31]);
        
    
        and(andpr29[32],b[28],a[32]);
        
    
        and(andpr29[33],b[28],a[33]);
        
    
        and(andpr29[34],b[28],a[34]);
        
    
        and(andpr29[35],b[28],a[35]);
        
    
        and(andpr29[36],b[28],a[36]);
        
    
        and(andpr29[37],b[28],a[37]);
        
    
        and(andpr29[38],b[28],a[38]);
        
    
        and(andpr29[39],b[28],a[39]);
        
    
        and(andpr29[40],b[28],a[40]);
        
    
        and(andpr29[41],b[28],a[41]);
        
    
        and(andpr29[42],b[28],a[42]);
        
    
        and(andpr29[43],b[28],a[43]);
        
    
        and(andpr29[44],b[28],a[44]);
        
    
        and(andpr29[45],b[28],a[45]);
        
    
        and(andpr29[46],b[28],a[46]);
        
    
        and(andpr29[47],b[28],a[47]);
        
    
        and(andpr29[48],b[28],a[48]);
        
    
        and(andpr29[49],b[28],a[49]);
        
    
        and(andpr29[50],b[28],a[50]);
        
    
        and(andpr29[51],b[28],a[51]);
        
    
        and(andpr29[52],b[28],a[52]);
        
    
        and(andpr29[53],b[28],a[53]);
        
    
        and(andpr29[54],b[28],a[54]);
        
    
        and(andpr29[55],b[28],a[55]);
        
    
        and(andpr29[56],b[28],a[56]);
        
    
        and(andpr29[57],b[28],a[57]);
        
    
        and(andpr29[58],b[28],a[58]);
        
    
        and(andpr29[59],b[28],a[59]);
        
    
        and(andpr29[60],b[28],a[60]);
        
    
        and(andpr29[61],b[28],a[61]);
        
    
        and(andpr29[62],b[28],a[62]);
        
    
        and(andpr29[63],b[28],a[63]);
        
    
    not(si[28],andpr29[63]);

    
        and(andpr30[0],b[29],a[0]);
        
    
        and(andpr30[1],b[29],a[1]);
        
    
        and(andpr30[2],b[29],a[2]);
        
    
        and(andpr30[3],b[29],a[3]);
        
    
        and(andpr30[4],b[29],a[4]);
        
    
        and(andpr30[5],b[29],a[5]);
        
    
        and(andpr30[6],b[29],a[6]);
        
    
        and(andpr30[7],b[29],a[7]);
        
    
        and(andpr30[8],b[29],a[8]);
        
    
        and(andpr30[9],b[29],a[9]);
        
    
        and(andpr30[10],b[29],a[10]);
        
    
        and(andpr30[11],b[29],a[11]);
        
    
        and(andpr30[12],b[29],a[12]);
        
    
        and(andpr30[13],b[29],a[13]);
        
    
        and(andpr30[14],b[29],a[14]);
        
    
        and(andpr30[15],b[29],a[15]);
        
    
        and(andpr30[16],b[29],a[16]);
        
    
        and(andpr30[17],b[29],a[17]);
        
    
        and(andpr30[18],b[29],a[18]);
        
    
        and(andpr30[19],b[29],a[19]);
        
    
        and(andpr30[20],b[29],a[20]);
        
    
        and(andpr30[21],b[29],a[21]);
        
    
        and(andpr30[22],b[29],a[22]);
        
    
        and(andpr30[23],b[29],a[23]);
        
    
        and(andpr30[24],b[29],a[24]);
        
    
        and(andpr30[25],b[29],a[25]);
        
    
        and(andpr30[26],b[29],a[26]);
        
    
        and(andpr30[27],b[29],a[27]);
        
    
        and(andpr30[28],b[29],a[28]);
        
    
        and(andpr30[29],b[29],a[29]);
        
    
        and(andpr30[30],b[29],a[30]);
        
    
        and(andpr30[31],b[29],a[31]);
        
    
        and(andpr30[32],b[29],a[32]);
        
    
        and(andpr30[33],b[29],a[33]);
        
    
        and(andpr30[34],b[29],a[34]);
        
    
        and(andpr30[35],b[29],a[35]);
        
    
        and(andpr30[36],b[29],a[36]);
        
    
        and(andpr30[37],b[29],a[37]);
        
    
        and(andpr30[38],b[29],a[38]);
        
    
        and(andpr30[39],b[29],a[39]);
        
    
        and(andpr30[40],b[29],a[40]);
        
    
        and(andpr30[41],b[29],a[41]);
        
    
        and(andpr30[42],b[29],a[42]);
        
    
        and(andpr30[43],b[29],a[43]);
        
    
        and(andpr30[44],b[29],a[44]);
        
    
        and(andpr30[45],b[29],a[45]);
        
    
        and(andpr30[46],b[29],a[46]);
        
    
        and(andpr30[47],b[29],a[47]);
        
    
        and(andpr30[48],b[29],a[48]);
        
    
        and(andpr30[49],b[29],a[49]);
        
    
        and(andpr30[50],b[29],a[50]);
        
    
        and(andpr30[51],b[29],a[51]);
        
    
        and(andpr30[52],b[29],a[52]);
        
    
        and(andpr30[53],b[29],a[53]);
        
    
        and(andpr30[54],b[29],a[54]);
        
    
        and(andpr30[55],b[29],a[55]);
        
    
        and(andpr30[56],b[29],a[56]);
        
    
        and(andpr30[57],b[29],a[57]);
        
    
        and(andpr30[58],b[29],a[58]);
        
    
        and(andpr30[59],b[29],a[59]);
        
    
        and(andpr30[60],b[29],a[60]);
        
    
        and(andpr30[61],b[29],a[61]);
        
    
        and(andpr30[62],b[29],a[62]);
        
    
        and(andpr30[63],b[29],a[63]);
        
    
    not(si[29],andpr30[63]);

    
        and(andpr31[0],b[30],a[0]);
        
    
        and(andpr31[1],b[30],a[1]);
        
    
        and(andpr31[2],b[30],a[2]);
        
    
        and(andpr31[3],b[30],a[3]);
        
    
        and(andpr31[4],b[30],a[4]);
        
    
        and(andpr31[5],b[30],a[5]);
        
    
        and(andpr31[6],b[30],a[6]);
        
    
        and(andpr31[7],b[30],a[7]);
        
    
        and(andpr31[8],b[30],a[8]);
        
    
        and(andpr31[9],b[30],a[9]);
        
    
        and(andpr31[10],b[30],a[10]);
        
    
        and(andpr31[11],b[30],a[11]);
        
    
        and(andpr31[12],b[30],a[12]);
        
    
        and(andpr31[13],b[30],a[13]);
        
    
        and(andpr31[14],b[30],a[14]);
        
    
        and(andpr31[15],b[30],a[15]);
        
    
        and(andpr31[16],b[30],a[16]);
        
    
        and(andpr31[17],b[30],a[17]);
        
    
        and(andpr31[18],b[30],a[18]);
        
    
        and(andpr31[19],b[30],a[19]);
        
    
        and(andpr31[20],b[30],a[20]);
        
    
        and(andpr31[21],b[30],a[21]);
        
    
        and(andpr31[22],b[30],a[22]);
        
    
        and(andpr31[23],b[30],a[23]);
        
    
        and(andpr31[24],b[30],a[24]);
        
    
        and(andpr31[25],b[30],a[25]);
        
    
        and(andpr31[26],b[30],a[26]);
        
    
        and(andpr31[27],b[30],a[27]);
        
    
        and(andpr31[28],b[30],a[28]);
        
    
        and(andpr31[29],b[30],a[29]);
        
    
        and(andpr31[30],b[30],a[30]);
        
    
        and(andpr31[31],b[30],a[31]);
        
    
        and(andpr31[32],b[30],a[32]);
        
    
        and(andpr31[33],b[30],a[33]);
        
    
        and(andpr31[34],b[30],a[34]);
        
    
        and(andpr31[35],b[30],a[35]);
        
    
        and(andpr31[36],b[30],a[36]);
        
    
        and(andpr31[37],b[30],a[37]);
        
    
        and(andpr31[38],b[30],a[38]);
        
    
        and(andpr31[39],b[30],a[39]);
        
    
        and(andpr31[40],b[30],a[40]);
        
    
        and(andpr31[41],b[30],a[41]);
        
    
        and(andpr31[42],b[30],a[42]);
        
    
        and(andpr31[43],b[30],a[43]);
        
    
        and(andpr31[44],b[30],a[44]);
        
    
        and(andpr31[45],b[30],a[45]);
        
    
        and(andpr31[46],b[30],a[46]);
        
    
        and(andpr31[47],b[30],a[47]);
        
    
        and(andpr31[48],b[30],a[48]);
        
    
        and(andpr31[49],b[30],a[49]);
        
    
        and(andpr31[50],b[30],a[50]);
        
    
        and(andpr31[51],b[30],a[51]);
        
    
        and(andpr31[52],b[30],a[52]);
        
    
        and(andpr31[53],b[30],a[53]);
        
    
        and(andpr31[54],b[30],a[54]);
        
    
        and(andpr31[55],b[30],a[55]);
        
    
        and(andpr31[56],b[30],a[56]);
        
    
        and(andpr31[57],b[30],a[57]);
        
    
        and(andpr31[58],b[30],a[58]);
        
    
        and(andpr31[59],b[30],a[59]);
        
    
        and(andpr31[60],b[30],a[60]);
        
    
        and(andpr31[61],b[30],a[61]);
        
    
        and(andpr31[62],b[30],a[62]);
        
    
        and(andpr31[63],b[30],a[63]);
        
    
    not(si[30],andpr31[63]);

    
        and(andpr32[0],b[31],a[0]);
        
    
        and(andpr32[1],b[31],a[1]);
        
    
        and(andpr32[2],b[31],a[2]);
        
    
        and(andpr32[3],b[31],a[3]);
        
    
        and(andpr32[4],b[31],a[4]);
        
    
        and(andpr32[5],b[31],a[5]);
        
    
        and(andpr32[6],b[31],a[6]);
        
    
        and(andpr32[7],b[31],a[7]);
        
    
        and(andpr32[8],b[31],a[8]);
        
    
        and(andpr32[9],b[31],a[9]);
        
    
        and(andpr32[10],b[31],a[10]);
        
    
        and(andpr32[11],b[31],a[11]);
        
    
        and(andpr32[12],b[31],a[12]);
        
    
        and(andpr32[13],b[31],a[13]);
        
    
        and(andpr32[14],b[31],a[14]);
        
    
        and(andpr32[15],b[31],a[15]);
        
    
        and(andpr32[16],b[31],a[16]);
        
    
        and(andpr32[17],b[31],a[17]);
        
    
        and(andpr32[18],b[31],a[18]);
        
    
        and(andpr32[19],b[31],a[19]);
        
    
        and(andpr32[20],b[31],a[20]);
        
    
        and(andpr32[21],b[31],a[21]);
        
    
        and(andpr32[22],b[31],a[22]);
        
    
        and(andpr32[23],b[31],a[23]);
        
    
        and(andpr32[24],b[31],a[24]);
        
    
        and(andpr32[25],b[31],a[25]);
        
    
        and(andpr32[26],b[31],a[26]);
        
    
        and(andpr32[27],b[31],a[27]);
        
    
        and(andpr32[28],b[31],a[28]);
        
    
        and(andpr32[29],b[31],a[29]);
        
    
        and(andpr32[30],b[31],a[30]);
        
    
        and(andpr32[31],b[31],a[31]);
        
    
        and(andpr32[32],b[31],a[32]);
        
    
        and(andpr32[33],b[31],a[33]);
        
    
        and(andpr32[34],b[31],a[34]);
        
    
        and(andpr32[35],b[31],a[35]);
        
    
        and(andpr32[36],b[31],a[36]);
        
    
        and(andpr32[37],b[31],a[37]);
        
    
        and(andpr32[38],b[31],a[38]);
        
    
        and(andpr32[39],b[31],a[39]);
        
    
        and(andpr32[40],b[31],a[40]);
        
    
        and(andpr32[41],b[31],a[41]);
        
    
        and(andpr32[42],b[31],a[42]);
        
    
        and(andpr32[43],b[31],a[43]);
        
    
        and(andpr32[44],b[31],a[44]);
        
    
        and(andpr32[45],b[31],a[45]);
        
    
        and(andpr32[46],b[31],a[46]);
        
    
        and(andpr32[47],b[31],a[47]);
        
    
        and(andpr32[48],b[31],a[48]);
        
    
        and(andpr32[49],b[31],a[49]);
        
    
        and(andpr32[50],b[31],a[50]);
        
    
        and(andpr32[51],b[31],a[51]);
        
    
        and(andpr32[52],b[31],a[52]);
        
    
        and(andpr32[53],b[31],a[53]);
        
    
        and(andpr32[54],b[31],a[54]);
        
    
        and(andpr32[55],b[31],a[55]);
        
    
        and(andpr32[56],b[31],a[56]);
        
    
        and(andpr32[57],b[31],a[57]);
        
    
        and(andpr32[58],b[31],a[58]);
        
    
        and(andpr32[59],b[31],a[59]);
        
    
        and(andpr32[60],b[31],a[60]);
        
    
        and(andpr32[61],b[31],a[61]);
        
    
        and(andpr32[62],b[31],a[62]);
        
    
        and(andpr32[63],b[31],a[63]);
        
    
    not(si[31],andpr32[63]);

    
        and(andpr33[0],b[32],a[0]);
        
    
        and(andpr33[1],b[32],a[1]);
        
    
        and(andpr33[2],b[32],a[2]);
        
    
        and(andpr33[3],b[32],a[3]);
        
    
        and(andpr33[4],b[32],a[4]);
        
    
        and(andpr33[5],b[32],a[5]);
        
    
        and(andpr33[6],b[32],a[6]);
        
    
        and(andpr33[7],b[32],a[7]);
        
    
        and(andpr33[8],b[32],a[8]);
        
    
        and(andpr33[9],b[32],a[9]);
        
    
        and(andpr33[10],b[32],a[10]);
        
    
        and(andpr33[11],b[32],a[11]);
        
    
        and(andpr33[12],b[32],a[12]);
        
    
        and(andpr33[13],b[32],a[13]);
        
    
        and(andpr33[14],b[32],a[14]);
        
    
        and(andpr33[15],b[32],a[15]);
        
    
        and(andpr33[16],b[32],a[16]);
        
    
        and(andpr33[17],b[32],a[17]);
        
    
        and(andpr33[18],b[32],a[18]);
        
    
        and(andpr33[19],b[32],a[19]);
        
    
        and(andpr33[20],b[32],a[20]);
        
    
        and(andpr33[21],b[32],a[21]);
        
    
        and(andpr33[22],b[32],a[22]);
        
    
        and(andpr33[23],b[32],a[23]);
        
    
        and(andpr33[24],b[32],a[24]);
        
    
        and(andpr33[25],b[32],a[25]);
        
    
        and(andpr33[26],b[32],a[26]);
        
    
        and(andpr33[27],b[32],a[27]);
        
    
        and(andpr33[28],b[32],a[28]);
        
    
        and(andpr33[29],b[32],a[29]);
        
    
        and(andpr33[30],b[32],a[30]);
        
    
        and(andpr33[31],b[32],a[31]);
        
    
        and(andpr33[32],b[32],a[32]);
        
    
        and(andpr33[33],b[32],a[33]);
        
    
        and(andpr33[34],b[32],a[34]);
        
    
        and(andpr33[35],b[32],a[35]);
        
    
        and(andpr33[36],b[32],a[36]);
        
    
        and(andpr33[37],b[32],a[37]);
        
    
        and(andpr33[38],b[32],a[38]);
        
    
        and(andpr33[39],b[32],a[39]);
        
    
        and(andpr33[40],b[32],a[40]);
        
    
        and(andpr33[41],b[32],a[41]);
        
    
        and(andpr33[42],b[32],a[42]);
        
    
        and(andpr33[43],b[32],a[43]);
        
    
        and(andpr33[44],b[32],a[44]);
        
    
        and(andpr33[45],b[32],a[45]);
        
    
        and(andpr33[46],b[32],a[46]);
        
    
        and(andpr33[47],b[32],a[47]);
        
    
        and(andpr33[48],b[32],a[48]);
        
    
        and(andpr33[49],b[32],a[49]);
        
    
        and(andpr33[50],b[32],a[50]);
        
    
        and(andpr33[51],b[32],a[51]);
        
    
        and(andpr33[52],b[32],a[52]);
        
    
        and(andpr33[53],b[32],a[53]);
        
    
        and(andpr33[54],b[32],a[54]);
        
    
        and(andpr33[55],b[32],a[55]);
        
    
        and(andpr33[56],b[32],a[56]);
        
    
        and(andpr33[57],b[32],a[57]);
        
    
        and(andpr33[58],b[32],a[58]);
        
    
        and(andpr33[59],b[32],a[59]);
        
    
        and(andpr33[60],b[32],a[60]);
        
    
        and(andpr33[61],b[32],a[61]);
        
    
        and(andpr33[62],b[32],a[62]);
        
    
        and(andpr33[63],b[32],a[63]);
        
    
    not(si[32],andpr33[63]);

    
        and(andpr34[0],b[33],a[0]);
        
    
        and(andpr34[1],b[33],a[1]);
        
    
        and(andpr34[2],b[33],a[2]);
        
    
        and(andpr34[3],b[33],a[3]);
        
    
        and(andpr34[4],b[33],a[4]);
        
    
        and(andpr34[5],b[33],a[5]);
        
    
        and(andpr34[6],b[33],a[6]);
        
    
        and(andpr34[7],b[33],a[7]);
        
    
        and(andpr34[8],b[33],a[8]);
        
    
        and(andpr34[9],b[33],a[9]);
        
    
        and(andpr34[10],b[33],a[10]);
        
    
        and(andpr34[11],b[33],a[11]);
        
    
        and(andpr34[12],b[33],a[12]);
        
    
        and(andpr34[13],b[33],a[13]);
        
    
        and(andpr34[14],b[33],a[14]);
        
    
        and(andpr34[15],b[33],a[15]);
        
    
        and(andpr34[16],b[33],a[16]);
        
    
        and(andpr34[17],b[33],a[17]);
        
    
        and(andpr34[18],b[33],a[18]);
        
    
        and(andpr34[19],b[33],a[19]);
        
    
        and(andpr34[20],b[33],a[20]);
        
    
        and(andpr34[21],b[33],a[21]);
        
    
        and(andpr34[22],b[33],a[22]);
        
    
        and(andpr34[23],b[33],a[23]);
        
    
        and(andpr34[24],b[33],a[24]);
        
    
        and(andpr34[25],b[33],a[25]);
        
    
        and(andpr34[26],b[33],a[26]);
        
    
        and(andpr34[27],b[33],a[27]);
        
    
        and(andpr34[28],b[33],a[28]);
        
    
        and(andpr34[29],b[33],a[29]);
        
    
        and(andpr34[30],b[33],a[30]);
        
    
        and(andpr34[31],b[33],a[31]);
        
    
        and(andpr34[32],b[33],a[32]);
        
    
        and(andpr34[33],b[33],a[33]);
        
    
        and(andpr34[34],b[33],a[34]);
        
    
        and(andpr34[35],b[33],a[35]);
        
    
        and(andpr34[36],b[33],a[36]);
        
    
        and(andpr34[37],b[33],a[37]);
        
    
        and(andpr34[38],b[33],a[38]);
        
    
        and(andpr34[39],b[33],a[39]);
        
    
        and(andpr34[40],b[33],a[40]);
        
    
        and(andpr34[41],b[33],a[41]);
        
    
        and(andpr34[42],b[33],a[42]);
        
    
        and(andpr34[43],b[33],a[43]);
        
    
        and(andpr34[44],b[33],a[44]);
        
    
        and(andpr34[45],b[33],a[45]);
        
    
        and(andpr34[46],b[33],a[46]);
        
    
        and(andpr34[47],b[33],a[47]);
        
    
        and(andpr34[48],b[33],a[48]);
        
    
        and(andpr34[49],b[33],a[49]);
        
    
        and(andpr34[50],b[33],a[50]);
        
    
        and(andpr34[51],b[33],a[51]);
        
    
        and(andpr34[52],b[33],a[52]);
        
    
        and(andpr34[53],b[33],a[53]);
        
    
        and(andpr34[54],b[33],a[54]);
        
    
        and(andpr34[55],b[33],a[55]);
        
    
        and(andpr34[56],b[33],a[56]);
        
    
        and(andpr34[57],b[33],a[57]);
        
    
        and(andpr34[58],b[33],a[58]);
        
    
        and(andpr34[59],b[33],a[59]);
        
    
        and(andpr34[60],b[33],a[60]);
        
    
        and(andpr34[61],b[33],a[61]);
        
    
        and(andpr34[62],b[33],a[62]);
        
    
        and(andpr34[63],b[33],a[63]);
        
    
    not(si[33],andpr34[63]);

    
        and(andpr35[0],b[34],a[0]);
        
    
        and(andpr35[1],b[34],a[1]);
        
    
        and(andpr35[2],b[34],a[2]);
        
    
        and(andpr35[3],b[34],a[3]);
        
    
        and(andpr35[4],b[34],a[4]);
        
    
        and(andpr35[5],b[34],a[5]);
        
    
        and(andpr35[6],b[34],a[6]);
        
    
        and(andpr35[7],b[34],a[7]);
        
    
        and(andpr35[8],b[34],a[8]);
        
    
        and(andpr35[9],b[34],a[9]);
        
    
        and(andpr35[10],b[34],a[10]);
        
    
        and(andpr35[11],b[34],a[11]);
        
    
        and(andpr35[12],b[34],a[12]);
        
    
        and(andpr35[13],b[34],a[13]);
        
    
        and(andpr35[14],b[34],a[14]);
        
    
        and(andpr35[15],b[34],a[15]);
        
    
        and(andpr35[16],b[34],a[16]);
        
    
        and(andpr35[17],b[34],a[17]);
        
    
        and(andpr35[18],b[34],a[18]);
        
    
        and(andpr35[19],b[34],a[19]);
        
    
        and(andpr35[20],b[34],a[20]);
        
    
        and(andpr35[21],b[34],a[21]);
        
    
        and(andpr35[22],b[34],a[22]);
        
    
        and(andpr35[23],b[34],a[23]);
        
    
        and(andpr35[24],b[34],a[24]);
        
    
        and(andpr35[25],b[34],a[25]);
        
    
        and(andpr35[26],b[34],a[26]);
        
    
        and(andpr35[27],b[34],a[27]);
        
    
        and(andpr35[28],b[34],a[28]);
        
    
        and(andpr35[29],b[34],a[29]);
        
    
        and(andpr35[30],b[34],a[30]);
        
    
        and(andpr35[31],b[34],a[31]);
        
    
        and(andpr35[32],b[34],a[32]);
        
    
        and(andpr35[33],b[34],a[33]);
        
    
        and(andpr35[34],b[34],a[34]);
        
    
        and(andpr35[35],b[34],a[35]);
        
    
        and(andpr35[36],b[34],a[36]);
        
    
        and(andpr35[37],b[34],a[37]);
        
    
        and(andpr35[38],b[34],a[38]);
        
    
        and(andpr35[39],b[34],a[39]);
        
    
        and(andpr35[40],b[34],a[40]);
        
    
        and(andpr35[41],b[34],a[41]);
        
    
        and(andpr35[42],b[34],a[42]);
        
    
        and(andpr35[43],b[34],a[43]);
        
    
        and(andpr35[44],b[34],a[44]);
        
    
        and(andpr35[45],b[34],a[45]);
        
    
        and(andpr35[46],b[34],a[46]);
        
    
        and(andpr35[47],b[34],a[47]);
        
    
        and(andpr35[48],b[34],a[48]);
        
    
        and(andpr35[49],b[34],a[49]);
        
    
        and(andpr35[50],b[34],a[50]);
        
    
        and(andpr35[51],b[34],a[51]);
        
    
        and(andpr35[52],b[34],a[52]);
        
    
        and(andpr35[53],b[34],a[53]);
        
    
        and(andpr35[54],b[34],a[54]);
        
    
        and(andpr35[55],b[34],a[55]);
        
    
        and(andpr35[56],b[34],a[56]);
        
    
        and(andpr35[57],b[34],a[57]);
        
    
        and(andpr35[58],b[34],a[58]);
        
    
        and(andpr35[59],b[34],a[59]);
        
    
        and(andpr35[60],b[34],a[60]);
        
    
        and(andpr35[61],b[34],a[61]);
        
    
        and(andpr35[62],b[34],a[62]);
        
    
        and(andpr35[63],b[34],a[63]);
        
    
    not(si[34],andpr35[63]);

    
        and(andpr36[0],b[35],a[0]);
        
    
        and(andpr36[1],b[35],a[1]);
        
    
        and(andpr36[2],b[35],a[2]);
        
    
        and(andpr36[3],b[35],a[3]);
        
    
        and(andpr36[4],b[35],a[4]);
        
    
        and(andpr36[5],b[35],a[5]);
        
    
        and(andpr36[6],b[35],a[6]);
        
    
        and(andpr36[7],b[35],a[7]);
        
    
        and(andpr36[8],b[35],a[8]);
        
    
        and(andpr36[9],b[35],a[9]);
        
    
        and(andpr36[10],b[35],a[10]);
        
    
        and(andpr36[11],b[35],a[11]);
        
    
        and(andpr36[12],b[35],a[12]);
        
    
        and(andpr36[13],b[35],a[13]);
        
    
        and(andpr36[14],b[35],a[14]);
        
    
        and(andpr36[15],b[35],a[15]);
        
    
        and(andpr36[16],b[35],a[16]);
        
    
        and(andpr36[17],b[35],a[17]);
        
    
        and(andpr36[18],b[35],a[18]);
        
    
        and(andpr36[19],b[35],a[19]);
        
    
        and(andpr36[20],b[35],a[20]);
        
    
        and(andpr36[21],b[35],a[21]);
        
    
        and(andpr36[22],b[35],a[22]);
        
    
        and(andpr36[23],b[35],a[23]);
        
    
        and(andpr36[24],b[35],a[24]);
        
    
        and(andpr36[25],b[35],a[25]);
        
    
        and(andpr36[26],b[35],a[26]);
        
    
        and(andpr36[27],b[35],a[27]);
        
    
        and(andpr36[28],b[35],a[28]);
        
    
        and(andpr36[29],b[35],a[29]);
        
    
        and(andpr36[30],b[35],a[30]);
        
    
        and(andpr36[31],b[35],a[31]);
        
    
        and(andpr36[32],b[35],a[32]);
        
    
        and(andpr36[33],b[35],a[33]);
        
    
        and(andpr36[34],b[35],a[34]);
        
    
        and(andpr36[35],b[35],a[35]);
        
    
        and(andpr36[36],b[35],a[36]);
        
    
        and(andpr36[37],b[35],a[37]);
        
    
        and(andpr36[38],b[35],a[38]);
        
    
        and(andpr36[39],b[35],a[39]);
        
    
        and(andpr36[40],b[35],a[40]);
        
    
        and(andpr36[41],b[35],a[41]);
        
    
        and(andpr36[42],b[35],a[42]);
        
    
        and(andpr36[43],b[35],a[43]);
        
    
        and(andpr36[44],b[35],a[44]);
        
    
        and(andpr36[45],b[35],a[45]);
        
    
        and(andpr36[46],b[35],a[46]);
        
    
        and(andpr36[47],b[35],a[47]);
        
    
        and(andpr36[48],b[35],a[48]);
        
    
        and(andpr36[49],b[35],a[49]);
        
    
        and(andpr36[50],b[35],a[50]);
        
    
        and(andpr36[51],b[35],a[51]);
        
    
        and(andpr36[52],b[35],a[52]);
        
    
        and(andpr36[53],b[35],a[53]);
        
    
        and(andpr36[54],b[35],a[54]);
        
    
        and(andpr36[55],b[35],a[55]);
        
    
        and(andpr36[56],b[35],a[56]);
        
    
        and(andpr36[57],b[35],a[57]);
        
    
        and(andpr36[58],b[35],a[58]);
        
    
        and(andpr36[59],b[35],a[59]);
        
    
        and(andpr36[60],b[35],a[60]);
        
    
        and(andpr36[61],b[35],a[61]);
        
    
        and(andpr36[62],b[35],a[62]);
        
    
        and(andpr36[63],b[35],a[63]);
        
    
    not(si[35],andpr36[63]);

    
        and(andpr37[0],b[36],a[0]);
        
    
        and(andpr37[1],b[36],a[1]);
        
    
        and(andpr37[2],b[36],a[2]);
        
    
        and(andpr37[3],b[36],a[3]);
        
    
        and(andpr37[4],b[36],a[4]);
        
    
        and(andpr37[5],b[36],a[5]);
        
    
        and(andpr37[6],b[36],a[6]);
        
    
        and(andpr37[7],b[36],a[7]);
        
    
        and(andpr37[8],b[36],a[8]);
        
    
        and(andpr37[9],b[36],a[9]);
        
    
        and(andpr37[10],b[36],a[10]);
        
    
        and(andpr37[11],b[36],a[11]);
        
    
        and(andpr37[12],b[36],a[12]);
        
    
        and(andpr37[13],b[36],a[13]);
        
    
        and(andpr37[14],b[36],a[14]);
        
    
        and(andpr37[15],b[36],a[15]);
        
    
        and(andpr37[16],b[36],a[16]);
        
    
        and(andpr37[17],b[36],a[17]);
        
    
        and(andpr37[18],b[36],a[18]);
        
    
        and(andpr37[19],b[36],a[19]);
        
    
        and(andpr37[20],b[36],a[20]);
        
    
        and(andpr37[21],b[36],a[21]);
        
    
        and(andpr37[22],b[36],a[22]);
        
    
        and(andpr37[23],b[36],a[23]);
        
    
        and(andpr37[24],b[36],a[24]);
        
    
        and(andpr37[25],b[36],a[25]);
        
    
        and(andpr37[26],b[36],a[26]);
        
    
        and(andpr37[27],b[36],a[27]);
        
    
        and(andpr37[28],b[36],a[28]);
        
    
        and(andpr37[29],b[36],a[29]);
        
    
        and(andpr37[30],b[36],a[30]);
        
    
        and(andpr37[31],b[36],a[31]);
        
    
        and(andpr37[32],b[36],a[32]);
        
    
        and(andpr37[33],b[36],a[33]);
        
    
        and(andpr37[34],b[36],a[34]);
        
    
        and(andpr37[35],b[36],a[35]);
        
    
        and(andpr37[36],b[36],a[36]);
        
    
        and(andpr37[37],b[36],a[37]);
        
    
        and(andpr37[38],b[36],a[38]);
        
    
        and(andpr37[39],b[36],a[39]);
        
    
        and(andpr37[40],b[36],a[40]);
        
    
        and(andpr37[41],b[36],a[41]);
        
    
        and(andpr37[42],b[36],a[42]);
        
    
        and(andpr37[43],b[36],a[43]);
        
    
        and(andpr37[44],b[36],a[44]);
        
    
        and(andpr37[45],b[36],a[45]);
        
    
        and(andpr37[46],b[36],a[46]);
        
    
        and(andpr37[47],b[36],a[47]);
        
    
        and(andpr37[48],b[36],a[48]);
        
    
        and(andpr37[49],b[36],a[49]);
        
    
        and(andpr37[50],b[36],a[50]);
        
    
        and(andpr37[51],b[36],a[51]);
        
    
        and(andpr37[52],b[36],a[52]);
        
    
        and(andpr37[53],b[36],a[53]);
        
    
        and(andpr37[54],b[36],a[54]);
        
    
        and(andpr37[55],b[36],a[55]);
        
    
        and(andpr37[56],b[36],a[56]);
        
    
        and(andpr37[57],b[36],a[57]);
        
    
        and(andpr37[58],b[36],a[58]);
        
    
        and(andpr37[59],b[36],a[59]);
        
    
        and(andpr37[60],b[36],a[60]);
        
    
        and(andpr37[61],b[36],a[61]);
        
    
        and(andpr37[62],b[36],a[62]);
        
    
        and(andpr37[63],b[36],a[63]);
        
    
    not(si[36],andpr37[63]);

    
        and(andpr38[0],b[37],a[0]);
        
    
        and(andpr38[1],b[37],a[1]);
        
    
        and(andpr38[2],b[37],a[2]);
        
    
        and(andpr38[3],b[37],a[3]);
        
    
        and(andpr38[4],b[37],a[4]);
        
    
        and(andpr38[5],b[37],a[5]);
        
    
        and(andpr38[6],b[37],a[6]);
        
    
        and(andpr38[7],b[37],a[7]);
        
    
        and(andpr38[8],b[37],a[8]);
        
    
        and(andpr38[9],b[37],a[9]);
        
    
        and(andpr38[10],b[37],a[10]);
        
    
        and(andpr38[11],b[37],a[11]);
        
    
        and(andpr38[12],b[37],a[12]);
        
    
        and(andpr38[13],b[37],a[13]);
        
    
        and(andpr38[14],b[37],a[14]);
        
    
        and(andpr38[15],b[37],a[15]);
        
    
        and(andpr38[16],b[37],a[16]);
        
    
        and(andpr38[17],b[37],a[17]);
        
    
        and(andpr38[18],b[37],a[18]);
        
    
        and(andpr38[19],b[37],a[19]);
        
    
        and(andpr38[20],b[37],a[20]);
        
    
        and(andpr38[21],b[37],a[21]);
        
    
        and(andpr38[22],b[37],a[22]);
        
    
        and(andpr38[23],b[37],a[23]);
        
    
        and(andpr38[24],b[37],a[24]);
        
    
        and(andpr38[25],b[37],a[25]);
        
    
        and(andpr38[26],b[37],a[26]);
        
    
        and(andpr38[27],b[37],a[27]);
        
    
        and(andpr38[28],b[37],a[28]);
        
    
        and(andpr38[29],b[37],a[29]);
        
    
        and(andpr38[30],b[37],a[30]);
        
    
        and(andpr38[31],b[37],a[31]);
        
    
        and(andpr38[32],b[37],a[32]);
        
    
        and(andpr38[33],b[37],a[33]);
        
    
        and(andpr38[34],b[37],a[34]);
        
    
        and(andpr38[35],b[37],a[35]);
        
    
        and(andpr38[36],b[37],a[36]);
        
    
        and(andpr38[37],b[37],a[37]);
        
    
        and(andpr38[38],b[37],a[38]);
        
    
        and(andpr38[39],b[37],a[39]);
        
    
        and(andpr38[40],b[37],a[40]);
        
    
        and(andpr38[41],b[37],a[41]);
        
    
        and(andpr38[42],b[37],a[42]);
        
    
        and(andpr38[43],b[37],a[43]);
        
    
        and(andpr38[44],b[37],a[44]);
        
    
        and(andpr38[45],b[37],a[45]);
        
    
        and(andpr38[46],b[37],a[46]);
        
    
        and(andpr38[47],b[37],a[47]);
        
    
        and(andpr38[48],b[37],a[48]);
        
    
        and(andpr38[49],b[37],a[49]);
        
    
        and(andpr38[50],b[37],a[50]);
        
    
        and(andpr38[51],b[37],a[51]);
        
    
        and(andpr38[52],b[37],a[52]);
        
    
        and(andpr38[53],b[37],a[53]);
        
    
        and(andpr38[54],b[37],a[54]);
        
    
        and(andpr38[55],b[37],a[55]);
        
    
        and(andpr38[56],b[37],a[56]);
        
    
        and(andpr38[57],b[37],a[57]);
        
    
        and(andpr38[58],b[37],a[58]);
        
    
        and(andpr38[59],b[37],a[59]);
        
    
        and(andpr38[60],b[37],a[60]);
        
    
        and(andpr38[61],b[37],a[61]);
        
    
        and(andpr38[62],b[37],a[62]);
        
    
        and(andpr38[63],b[37],a[63]);
        
    
    not(si[37],andpr38[63]);

    
        and(andpr39[0],b[38],a[0]);
        
    
        and(andpr39[1],b[38],a[1]);
        
    
        and(andpr39[2],b[38],a[2]);
        
    
        and(andpr39[3],b[38],a[3]);
        
    
        and(andpr39[4],b[38],a[4]);
        
    
        and(andpr39[5],b[38],a[5]);
        
    
        and(andpr39[6],b[38],a[6]);
        
    
        and(andpr39[7],b[38],a[7]);
        
    
        and(andpr39[8],b[38],a[8]);
        
    
        and(andpr39[9],b[38],a[9]);
        
    
        and(andpr39[10],b[38],a[10]);
        
    
        and(andpr39[11],b[38],a[11]);
        
    
        and(andpr39[12],b[38],a[12]);
        
    
        and(andpr39[13],b[38],a[13]);
        
    
        and(andpr39[14],b[38],a[14]);
        
    
        and(andpr39[15],b[38],a[15]);
        
    
        and(andpr39[16],b[38],a[16]);
        
    
        and(andpr39[17],b[38],a[17]);
        
    
        and(andpr39[18],b[38],a[18]);
        
    
        and(andpr39[19],b[38],a[19]);
        
    
        and(andpr39[20],b[38],a[20]);
        
    
        and(andpr39[21],b[38],a[21]);
        
    
        and(andpr39[22],b[38],a[22]);
        
    
        and(andpr39[23],b[38],a[23]);
        
    
        and(andpr39[24],b[38],a[24]);
        
    
        and(andpr39[25],b[38],a[25]);
        
    
        and(andpr39[26],b[38],a[26]);
        
    
        and(andpr39[27],b[38],a[27]);
        
    
        and(andpr39[28],b[38],a[28]);
        
    
        and(andpr39[29],b[38],a[29]);
        
    
        and(andpr39[30],b[38],a[30]);
        
    
        and(andpr39[31],b[38],a[31]);
        
    
        and(andpr39[32],b[38],a[32]);
        
    
        and(andpr39[33],b[38],a[33]);
        
    
        and(andpr39[34],b[38],a[34]);
        
    
        and(andpr39[35],b[38],a[35]);
        
    
        and(andpr39[36],b[38],a[36]);
        
    
        and(andpr39[37],b[38],a[37]);
        
    
        and(andpr39[38],b[38],a[38]);
        
    
        and(andpr39[39],b[38],a[39]);
        
    
        and(andpr39[40],b[38],a[40]);
        
    
        and(andpr39[41],b[38],a[41]);
        
    
        and(andpr39[42],b[38],a[42]);
        
    
        and(andpr39[43],b[38],a[43]);
        
    
        and(andpr39[44],b[38],a[44]);
        
    
        and(andpr39[45],b[38],a[45]);
        
    
        and(andpr39[46],b[38],a[46]);
        
    
        and(andpr39[47],b[38],a[47]);
        
    
        and(andpr39[48],b[38],a[48]);
        
    
        and(andpr39[49],b[38],a[49]);
        
    
        and(andpr39[50],b[38],a[50]);
        
    
        and(andpr39[51],b[38],a[51]);
        
    
        and(andpr39[52],b[38],a[52]);
        
    
        and(andpr39[53],b[38],a[53]);
        
    
        and(andpr39[54],b[38],a[54]);
        
    
        and(andpr39[55],b[38],a[55]);
        
    
        and(andpr39[56],b[38],a[56]);
        
    
        and(andpr39[57],b[38],a[57]);
        
    
        and(andpr39[58],b[38],a[58]);
        
    
        and(andpr39[59],b[38],a[59]);
        
    
        and(andpr39[60],b[38],a[60]);
        
    
        and(andpr39[61],b[38],a[61]);
        
    
        and(andpr39[62],b[38],a[62]);
        
    
        and(andpr39[63],b[38],a[63]);
        
    
    not(si[38],andpr39[63]);

    
        and(andpr40[0],b[39],a[0]);
        
    
        and(andpr40[1],b[39],a[1]);
        
    
        and(andpr40[2],b[39],a[2]);
        
    
        and(andpr40[3],b[39],a[3]);
        
    
        and(andpr40[4],b[39],a[4]);
        
    
        and(andpr40[5],b[39],a[5]);
        
    
        and(andpr40[6],b[39],a[6]);
        
    
        and(andpr40[7],b[39],a[7]);
        
    
        and(andpr40[8],b[39],a[8]);
        
    
        and(andpr40[9],b[39],a[9]);
        
    
        and(andpr40[10],b[39],a[10]);
        
    
        and(andpr40[11],b[39],a[11]);
        
    
        and(andpr40[12],b[39],a[12]);
        
    
        and(andpr40[13],b[39],a[13]);
        
    
        and(andpr40[14],b[39],a[14]);
        
    
        and(andpr40[15],b[39],a[15]);
        
    
        and(andpr40[16],b[39],a[16]);
        
    
        and(andpr40[17],b[39],a[17]);
        
    
        and(andpr40[18],b[39],a[18]);
        
    
        and(andpr40[19],b[39],a[19]);
        
    
        and(andpr40[20],b[39],a[20]);
        
    
        and(andpr40[21],b[39],a[21]);
        
    
        and(andpr40[22],b[39],a[22]);
        
    
        and(andpr40[23],b[39],a[23]);
        
    
        and(andpr40[24],b[39],a[24]);
        
    
        and(andpr40[25],b[39],a[25]);
        
    
        and(andpr40[26],b[39],a[26]);
        
    
        and(andpr40[27],b[39],a[27]);
        
    
        and(andpr40[28],b[39],a[28]);
        
    
        and(andpr40[29],b[39],a[29]);
        
    
        and(andpr40[30],b[39],a[30]);
        
    
        and(andpr40[31],b[39],a[31]);
        
    
        and(andpr40[32],b[39],a[32]);
        
    
        and(andpr40[33],b[39],a[33]);
        
    
        and(andpr40[34],b[39],a[34]);
        
    
        and(andpr40[35],b[39],a[35]);
        
    
        and(andpr40[36],b[39],a[36]);
        
    
        and(andpr40[37],b[39],a[37]);
        
    
        and(andpr40[38],b[39],a[38]);
        
    
        and(andpr40[39],b[39],a[39]);
        
    
        and(andpr40[40],b[39],a[40]);
        
    
        and(andpr40[41],b[39],a[41]);
        
    
        and(andpr40[42],b[39],a[42]);
        
    
        and(andpr40[43],b[39],a[43]);
        
    
        and(andpr40[44],b[39],a[44]);
        
    
        and(andpr40[45],b[39],a[45]);
        
    
        and(andpr40[46],b[39],a[46]);
        
    
        and(andpr40[47],b[39],a[47]);
        
    
        and(andpr40[48],b[39],a[48]);
        
    
        and(andpr40[49],b[39],a[49]);
        
    
        and(andpr40[50],b[39],a[50]);
        
    
        and(andpr40[51],b[39],a[51]);
        
    
        and(andpr40[52],b[39],a[52]);
        
    
        and(andpr40[53],b[39],a[53]);
        
    
        and(andpr40[54],b[39],a[54]);
        
    
        and(andpr40[55],b[39],a[55]);
        
    
        and(andpr40[56],b[39],a[56]);
        
    
        and(andpr40[57],b[39],a[57]);
        
    
        and(andpr40[58],b[39],a[58]);
        
    
        and(andpr40[59],b[39],a[59]);
        
    
        and(andpr40[60],b[39],a[60]);
        
    
        and(andpr40[61],b[39],a[61]);
        
    
        and(andpr40[62],b[39],a[62]);
        
    
        and(andpr40[63],b[39],a[63]);
        
    
    not(si[39],andpr40[63]);

    
        and(andpr41[0],b[40],a[0]);
        
    
        and(andpr41[1],b[40],a[1]);
        
    
        and(andpr41[2],b[40],a[2]);
        
    
        and(andpr41[3],b[40],a[3]);
        
    
        and(andpr41[4],b[40],a[4]);
        
    
        and(andpr41[5],b[40],a[5]);
        
    
        and(andpr41[6],b[40],a[6]);
        
    
        and(andpr41[7],b[40],a[7]);
        
    
        and(andpr41[8],b[40],a[8]);
        
    
        and(andpr41[9],b[40],a[9]);
        
    
        and(andpr41[10],b[40],a[10]);
        
    
        and(andpr41[11],b[40],a[11]);
        
    
        and(andpr41[12],b[40],a[12]);
        
    
        and(andpr41[13],b[40],a[13]);
        
    
        and(andpr41[14],b[40],a[14]);
        
    
        and(andpr41[15],b[40],a[15]);
        
    
        and(andpr41[16],b[40],a[16]);
        
    
        and(andpr41[17],b[40],a[17]);
        
    
        and(andpr41[18],b[40],a[18]);
        
    
        and(andpr41[19],b[40],a[19]);
        
    
        and(andpr41[20],b[40],a[20]);
        
    
        and(andpr41[21],b[40],a[21]);
        
    
        and(andpr41[22],b[40],a[22]);
        
    
        and(andpr41[23],b[40],a[23]);
        
    
        and(andpr41[24],b[40],a[24]);
        
    
        and(andpr41[25],b[40],a[25]);
        
    
        and(andpr41[26],b[40],a[26]);
        
    
        and(andpr41[27],b[40],a[27]);
        
    
        and(andpr41[28],b[40],a[28]);
        
    
        and(andpr41[29],b[40],a[29]);
        
    
        and(andpr41[30],b[40],a[30]);
        
    
        and(andpr41[31],b[40],a[31]);
        
    
        and(andpr41[32],b[40],a[32]);
        
    
        and(andpr41[33],b[40],a[33]);
        
    
        and(andpr41[34],b[40],a[34]);
        
    
        and(andpr41[35],b[40],a[35]);
        
    
        and(andpr41[36],b[40],a[36]);
        
    
        and(andpr41[37],b[40],a[37]);
        
    
        and(andpr41[38],b[40],a[38]);
        
    
        and(andpr41[39],b[40],a[39]);
        
    
        and(andpr41[40],b[40],a[40]);
        
    
        and(andpr41[41],b[40],a[41]);
        
    
        and(andpr41[42],b[40],a[42]);
        
    
        and(andpr41[43],b[40],a[43]);
        
    
        and(andpr41[44],b[40],a[44]);
        
    
        and(andpr41[45],b[40],a[45]);
        
    
        and(andpr41[46],b[40],a[46]);
        
    
        and(andpr41[47],b[40],a[47]);
        
    
        and(andpr41[48],b[40],a[48]);
        
    
        and(andpr41[49],b[40],a[49]);
        
    
        and(andpr41[50],b[40],a[50]);
        
    
        and(andpr41[51],b[40],a[51]);
        
    
        and(andpr41[52],b[40],a[52]);
        
    
        and(andpr41[53],b[40],a[53]);
        
    
        and(andpr41[54],b[40],a[54]);
        
    
        and(andpr41[55],b[40],a[55]);
        
    
        and(andpr41[56],b[40],a[56]);
        
    
        and(andpr41[57],b[40],a[57]);
        
    
        and(andpr41[58],b[40],a[58]);
        
    
        and(andpr41[59],b[40],a[59]);
        
    
        and(andpr41[60],b[40],a[60]);
        
    
        and(andpr41[61],b[40],a[61]);
        
    
        and(andpr41[62],b[40],a[62]);
        
    
        and(andpr41[63],b[40],a[63]);
        
    
    not(si[40],andpr41[63]);

    
        and(andpr42[0],b[41],a[0]);
        
    
        and(andpr42[1],b[41],a[1]);
        
    
        and(andpr42[2],b[41],a[2]);
        
    
        and(andpr42[3],b[41],a[3]);
        
    
        and(andpr42[4],b[41],a[4]);
        
    
        and(andpr42[5],b[41],a[5]);
        
    
        and(andpr42[6],b[41],a[6]);
        
    
        and(andpr42[7],b[41],a[7]);
        
    
        and(andpr42[8],b[41],a[8]);
        
    
        and(andpr42[9],b[41],a[9]);
        
    
        and(andpr42[10],b[41],a[10]);
        
    
        and(andpr42[11],b[41],a[11]);
        
    
        and(andpr42[12],b[41],a[12]);
        
    
        and(andpr42[13],b[41],a[13]);
        
    
        and(andpr42[14],b[41],a[14]);
        
    
        and(andpr42[15],b[41],a[15]);
        
    
        and(andpr42[16],b[41],a[16]);
        
    
        and(andpr42[17],b[41],a[17]);
        
    
        and(andpr42[18],b[41],a[18]);
        
    
        and(andpr42[19],b[41],a[19]);
        
    
        and(andpr42[20],b[41],a[20]);
        
    
        and(andpr42[21],b[41],a[21]);
        
    
        and(andpr42[22],b[41],a[22]);
        
    
        and(andpr42[23],b[41],a[23]);
        
    
        and(andpr42[24],b[41],a[24]);
        
    
        and(andpr42[25],b[41],a[25]);
        
    
        and(andpr42[26],b[41],a[26]);
        
    
        and(andpr42[27],b[41],a[27]);
        
    
        and(andpr42[28],b[41],a[28]);
        
    
        and(andpr42[29],b[41],a[29]);
        
    
        and(andpr42[30],b[41],a[30]);
        
    
        and(andpr42[31],b[41],a[31]);
        
    
        and(andpr42[32],b[41],a[32]);
        
    
        and(andpr42[33],b[41],a[33]);
        
    
        and(andpr42[34],b[41],a[34]);
        
    
        and(andpr42[35],b[41],a[35]);
        
    
        and(andpr42[36],b[41],a[36]);
        
    
        and(andpr42[37],b[41],a[37]);
        
    
        and(andpr42[38],b[41],a[38]);
        
    
        and(andpr42[39],b[41],a[39]);
        
    
        and(andpr42[40],b[41],a[40]);
        
    
        and(andpr42[41],b[41],a[41]);
        
    
        and(andpr42[42],b[41],a[42]);
        
    
        and(andpr42[43],b[41],a[43]);
        
    
        and(andpr42[44],b[41],a[44]);
        
    
        and(andpr42[45],b[41],a[45]);
        
    
        and(andpr42[46],b[41],a[46]);
        
    
        and(andpr42[47],b[41],a[47]);
        
    
        and(andpr42[48],b[41],a[48]);
        
    
        and(andpr42[49],b[41],a[49]);
        
    
        and(andpr42[50],b[41],a[50]);
        
    
        and(andpr42[51],b[41],a[51]);
        
    
        and(andpr42[52],b[41],a[52]);
        
    
        and(andpr42[53],b[41],a[53]);
        
    
        and(andpr42[54],b[41],a[54]);
        
    
        and(andpr42[55],b[41],a[55]);
        
    
        and(andpr42[56],b[41],a[56]);
        
    
        and(andpr42[57],b[41],a[57]);
        
    
        and(andpr42[58],b[41],a[58]);
        
    
        and(andpr42[59],b[41],a[59]);
        
    
        and(andpr42[60],b[41],a[60]);
        
    
        and(andpr42[61],b[41],a[61]);
        
    
        and(andpr42[62],b[41],a[62]);
        
    
        and(andpr42[63],b[41],a[63]);
        
    
    not(si[41],andpr42[63]);

    
        and(andpr43[0],b[42],a[0]);
        
    
        and(andpr43[1],b[42],a[1]);
        
    
        and(andpr43[2],b[42],a[2]);
        
    
        and(andpr43[3],b[42],a[3]);
        
    
        and(andpr43[4],b[42],a[4]);
        
    
        and(andpr43[5],b[42],a[5]);
        
    
        and(andpr43[6],b[42],a[6]);
        
    
        and(andpr43[7],b[42],a[7]);
        
    
        and(andpr43[8],b[42],a[8]);
        
    
        and(andpr43[9],b[42],a[9]);
        
    
        and(andpr43[10],b[42],a[10]);
        
    
        and(andpr43[11],b[42],a[11]);
        
    
        and(andpr43[12],b[42],a[12]);
        
    
        and(andpr43[13],b[42],a[13]);
        
    
        and(andpr43[14],b[42],a[14]);
        
    
        and(andpr43[15],b[42],a[15]);
        
    
        and(andpr43[16],b[42],a[16]);
        
    
        and(andpr43[17],b[42],a[17]);
        
    
        and(andpr43[18],b[42],a[18]);
        
    
        and(andpr43[19],b[42],a[19]);
        
    
        and(andpr43[20],b[42],a[20]);
        
    
        and(andpr43[21],b[42],a[21]);
        
    
        and(andpr43[22],b[42],a[22]);
        
    
        and(andpr43[23],b[42],a[23]);
        
    
        and(andpr43[24],b[42],a[24]);
        
    
        and(andpr43[25],b[42],a[25]);
        
    
        and(andpr43[26],b[42],a[26]);
        
    
        and(andpr43[27],b[42],a[27]);
        
    
        and(andpr43[28],b[42],a[28]);
        
    
        and(andpr43[29],b[42],a[29]);
        
    
        and(andpr43[30],b[42],a[30]);
        
    
        and(andpr43[31],b[42],a[31]);
        
    
        and(andpr43[32],b[42],a[32]);
        
    
        and(andpr43[33],b[42],a[33]);
        
    
        and(andpr43[34],b[42],a[34]);
        
    
        and(andpr43[35],b[42],a[35]);
        
    
        and(andpr43[36],b[42],a[36]);
        
    
        and(andpr43[37],b[42],a[37]);
        
    
        and(andpr43[38],b[42],a[38]);
        
    
        and(andpr43[39],b[42],a[39]);
        
    
        and(andpr43[40],b[42],a[40]);
        
    
        and(andpr43[41],b[42],a[41]);
        
    
        and(andpr43[42],b[42],a[42]);
        
    
        and(andpr43[43],b[42],a[43]);
        
    
        and(andpr43[44],b[42],a[44]);
        
    
        and(andpr43[45],b[42],a[45]);
        
    
        and(andpr43[46],b[42],a[46]);
        
    
        and(andpr43[47],b[42],a[47]);
        
    
        and(andpr43[48],b[42],a[48]);
        
    
        and(andpr43[49],b[42],a[49]);
        
    
        and(andpr43[50],b[42],a[50]);
        
    
        and(andpr43[51],b[42],a[51]);
        
    
        and(andpr43[52],b[42],a[52]);
        
    
        and(andpr43[53],b[42],a[53]);
        
    
        and(andpr43[54],b[42],a[54]);
        
    
        and(andpr43[55],b[42],a[55]);
        
    
        and(andpr43[56],b[42],a[56]);
        
    
        and(andpr43[57],b[42],a[57]);
        
    
        and(andpr43[58],b[42],a[58]);
        
    
        and(andpr43[59],b[42],a[59]);
        
    
        and(andpr43[60],b[42],a[60]);
        
    
        and(andpr43[61],b[42],a[61]);
        
    
        and(andpr43[62],b[42],a[62]);
        
    
        and(andpr43[63],b[42],a[63]);
        
    
    not(si[42],andpr43[63]);

    
        and(andpr44[0],b[43],a[0]);
        
    
        and(andpr44[1],b[43],a[1]);
        
    
        and(andpr44[2],b[43],a[2]);
        
    
        and(andpr44[3],b[43],a[3]);
        
    
        and(andpr44[4],b[43],a[4]);
        
    
        and(andpr44[5],b[43],a[5]);
        
    
        and(andpr44[6],b[43],a[6]);
        
    
        and(andpr44[7],b[43],a[7]);
        
    
        and(andpr44[8],b[43],a[8]);
        
    
        and(andpr44[9],b[43],a[9]);
        
    
        and(andpr44[10],b[43],a[10]);
        
    
        and(andpr44[11],b[43],a[11]);
        
    
        and(andpr44[12],b[43],a[12]);
        
    
        and(andpr44[13],b[43],a[13]);
        
    
        and(andpr44[14],b[43],a[14]);
        
    
        and(andpr44[15],b[43],a[15]);
        
    
        and(andpr44[16],b[43],a[16]);
        
    
        and(andpr44[17],b[43],a[17]);
        
    
        and(andpr44[18],b[43],a[18]);
        
    
        and(andpr44[19],b[43],a[19]);
        
    
        and(andpr44[20],b[43],a[20]);
        
    
        and(andpr44[21],b[43],a[21]);
        
    
        and(andpr44[22],b[43],a[22]);
        
    
        and(andpr44[23],b[43],a[23]);
        
    
        and(andpr44[24],b[43],a[24]);
        
    
        and(andpr44[25],b[43],a[25]);
        
    
        and(andpr44[26],b[43],a[26]);
        
    
        and(andpr44[27],b[43],a[27]);
        
    
        and(andpr44[28],b[43],a[28]);
        
    
        and(andpr44[29],b[43],a[29]);
        
    
        and(andpr44[30],b[43],a[30]);
        
    
        and(andpr44[31],b[43],a[31]);
        
    
        and(andpr44[32],b[43],a[32]);
        
    
        and(andpr44[33],b[43],a[33]);
        
    
        and(andpr44[34],b[43],a[34]);
        
    
        and(andpr44[35],b[43],a[35]);
        
    
        and(andpr44[36],b[43],a[36]);
        
    
        and(andpr44[37],b[43],a[37]);
        
    
        and(andpr44[38],b[43],a[38]);
        
    
        and(andpr44[39],b[43],a[39]);
        
    
        and(andpr44[40],b[43],a[40]);
        
    
        and(andpr44[41],b[43],a[41]);
        
    
        and(andpr44[42],b[43],a[42]);
        
    
        and(andpr44[43],b[43],a[43]);
        
    
        and(andpr44[44],b[43],a[44]);
        
    
        and(andpr44[45],b[43],a[45]);
        
    
        and(andpr44[46],b[43],a[46]);
        
    
        and(andpr44[47],b[43],a[47]);
        
    
        and(andpr44[48],b[43],a[48]);
        
    
        and(andpr44[49],b[43],a[49]);
        
    
        and(andpr44[50],b[43],a[50]);
        
    
        and(andpr44[51],b[43],a[51]);
        
    
        and(andpr44[52],b[43],a[52]);
        
    
        and(andpr44[53],b[43],a[53]);
        
    
        and(andpr44[54],b[43],a[54]);
        
    
        and(andpr44[55],b[43],a[55]);
        
    
        and(andpr44[56],b[43],a[56]);
        
    
        and(andpr44[57],b[43],a[57]);
        
    
        and(andpr44[58],b[43],a[58]);
        
    
        and(andpr44[59],b[43],a[59]);
        
    
        and(andpr44[60],b[43],a[60]);
        
    
        and(andpr44[61],b[43],a[61]);
        
    
        and(andpr44[62],b[43],a[62]);
        
    
        and(andpr44[63],b[43],a[63]);
        
    
    not(si[43],andpr44[63]);

    
        and(andpr45[0],b[44],a[0]);
        
    
        and(andpr45[1],b[44],a[1]);
        
    
        and(andpr45[2],b[44],a[2]);
        
    
        and(andpr45[3],b[44],a[3]);
        
    
        and(andpr45[4],b[44],a[4]);
        
    
        and(andpr45[5],b[44],a[5]);
        
    
        and(andpr45[6],b[44],a[6]);
        
    
        and(andpr45[7],b[44],a[7]);
        
    
        and(andpr45[8],b[44],a[8]);
        
    
        and(andpr45[9],b[44],a[9]);
        
    
        and(andpr45[10],b[44],a[10]);
        
    
        and(andpr45[11],b[44],a[11]);
        
    
        and(andpr45[12],b[44],a[12]);
        
    
        and(andpr45[13],b[44],a[13]);
        
    
        and(andpr45[14],b[44],a[14]);
        
    
        and(andpr45[15],b[44],a[15]);
        
    
        and(andpr45[16],b[44],a[16]);
        
    
        and(andpr45[17],b[44],a[17]);
        
    
        and(andpr45[18],b[44],a[18]);
        
    
        and(andpr45[19],b[44],a[19]);
        
    
        and(andpr45[20],b[44],a[20]);
        
    
        and(andpr45[21],b[44],a[21]);
        
    
        and(andpr45[22],b[44],a[22]);
        
    
        and(andpr45[23],b[44],a[23]);
        
    
        and(andpr45[24],b[44],a[24]);
        
    
        and(andpr45[25],b[44],a[25]);
        
    
        and(andpr45[26],b[44],a[26]);
        
    
        and(andpr45[27],b[44],a[27]);
        
    
        and(andpr45[28],b[44],a[28]);
        
    
        and(andpr45[29],b[44],a[29]);
        
    
        and(andpr45[30],b[44],a[30]);
        
    
        and(andpr45[31],b[44],a[31]);
        
    
        and(andpr45[32],b[44],a[32]);
        
    
        and(andpr45[33],b[44],a[33]);
        
    
        and(andpr45[34],b[44],a[34]);
        
    
        and(andpr45[35],b[44],a[35]);
        
    
        and(andpr45[36],b[44],a[36]);
        
    
        and(andpr45[37],b[44],a[37]);
        
    
        and(andpr45[38],b[44],a[38]);
        
    
        and(andpr45[39],b[44],a[39]);
        
    
        and(andpr45[40],b[44],a[40]);
        
    
        and(andpr45[41],b[44],a[41]);
        
    
        and(andpr45[42],b[44],a[42]);
        
    
        and(andpr45[43],b[44],a[43]);
        
    
        and(andpr45[44],b[44],a[44]);
        
    
        and(andpr45[45],b[44],a[45]);
        
    
        and(andpr45[46],b[44],a[46]);
        
    
        and(andpr45[47],b[44],a[47]);
        
    
        and(andpr45[48],b[44],a[48]);
        
    
        and(andpr45[49],b[44],a[49]);
        
    
        and(andpr45[50],b[44],a[50]);
        
    
        and(andpr45[51],b[44],a[51]);
        
    
        and(andpr45[52],b[44],a[52]);
        
    
        and(andpr45[53],b[44],a[53]);
        
    
        and(andpr45[54],b[44],a[54]);
        
    
        and(andpr45[55],b[44],a[55]);
        
    
        and(andpr45[56],b[44],a[56]);
        
    
        and(andpr45[57],b[44],a[57]);
        
    
        and(andpr45[58],b[44],a[58]);
        
    
        and(andpr45[59],b[44],a[59]);
        
    
        and(andpr45[60],b[44],a[60]);
        
    
        and(andpr45[61],b[44],a[61]);
        
    
        and(andpr45[62],b[44],a[62]);
        
    
        and(andpr45[63],b[44],a[63]);
        
    
    not(si[44],andpr45[63]);

    
        and(andpr46[0],b[45],a[0]);
        
    
        and(andpr46[1],b[45],a[1]);
        
    
        and(andpr46[2],b[45],a[2]);
        
    
        and(andpr46[3],b[45],a[3]);
        
    
        and(andpr46[4],b[45],a[4]);
        
    
        and(andpr46[5],b[45],a[5]);
        
    
        and(andpr46[6],b[45],a[6]);
        
    
        and(andpr46[7],b[45],a[7]);
        
    
        and(andpr46[8],b[45],a[8]);
        
    
        and(andpr46[9],b[45],a[9]);
        
    
        and(andpr46[10],b[45],a[10]);
        
    
        and(andpr46[11],b[45],a[11]);
        
    
        and(andpr46[12],b[45],a[12]);
        
    
        and(andpr46[13],b[45],a[13]);
        
    
        and(andpr46[14],b[45],a[14]);
        
    
        and(andpr46[15],b[45],a[15]);
        
    
        and(andpr46[16],b[45],a[16]);
        
    
        and(andpr46[17],b[45],a[17]);
        
    
        and(andpr46[18],b[45],a[18]);
        
    
        and(andpr46[19],b[45],a[19]);
        
    
        and(andpr46[20],b[45],a[20]);
        
    
        and(andpr46[21],b[45],a[21]);
        
    
        and(andpr46[22],b[45],a[22]);
        
    
        and(andpr46[23],b[45],a[23]);
        
    
        and(andpr46[24],b[45],a[24]);
        
    
        and(andpr46[25],b[45],a[25]);
        
    
        and(andpr46[26],b[45],a[26]);
        
    
        and(andpr46[27],b[45],a[27]);
        
    
        and(andpr46[28],b[45],a[28]);
        
    
        and(andpr46[29],b[45],a[29]);
        
    
        and(andpr46[30],b[45],a[30]);
        
    
        and(andpr46[31],b[45],a[31]);
        
    
        and(andpr46[32],b[45],a[32]);
        
    
        and(andpr46[33],b[45],a[33]);
        
    
        and(andpr46[34],b[45],a[34]);
        
    
        and(andpr46[35],b[45],a[35]);
        
    
        and(andpr46[36],b[45],a[36]);
        
    
        and(andpr46[37],b[45],a[37]);
        
    
        and(andpr46[38],b[45],a[38]);
        
    
        and(andpr46[39],b[45],a[39]);
        
    
        and(andpr46[40],b[45],a[40]);
        
    
        and(andpr46[41],b[45],a[41]);
        
    
        and(andpr46[42],b[45],a[42]);
        
    
        and(andpr46[43],b[45],a[43]);
        
    
        and(andpr46[44],b[45],a[44]);
        
    
        and(andpr46[45],b[45],a[45]);
        
    
        and(andpr46[46],b[45],a[46]);
        
    
        and(andpr46[47],b[45],a[47]);
        
    
        and(andpr46[48],b[45],a[48]);
        
    
        and(andpr46[49],b[45],a[49]);
        
    
        and(andpr46[50],b[45],a[50]);
        
    
        and(andpr46[51],b[45],a[51]);
        
    
        and(andpr46[52],b[45],a[52]);
        
    
        and(andpr46[53],b[45],a[53]);
        
    
        and(andpr46[54],b[45],a[54]);
        
    
        and(andpr46[55],b[45],a[55]);
        
    
        and(andpr46[56],b[45],a[56]);
        
    
        and(andpr46[57],b[45],a[57]);
        
    
        and(andpr46[58],b[45],a[58]);
        
    
        and(andpr46[59],b[45],a[59]);
        
    
        and(andpr46[60],b[45],a[60]);
        
    
        and(andpr46[61],b[45],a[61]);
        
    
        and(andpr46[62],b[45],a[62]);
        
    
        and(andpr46[63],b[45],a[63]);
        
    
    not(si[45],andpr46[63]);

    
        and(andpr47[0],b[46],a[0]);
        
    
        and(andpr47[1],b[46],a[1]);
        
    
        and(andpr47[2],b[46],a[2]);
        
    
        and(andpr47[3],b[46],a[3]);
        
    
        and(andpr47[4],b[46],a[4]);
        
    
        and(andpr47[5],b[46],a[5]);
        
    
        and(andpr47[6],b[46],a[6]);
        
    
        and(andpr47[7],b[46],a[7]);
        
    
        and(andpr47[8],b[46],a[8]);
        
    
        and(andpr47[9],b[46],a[9]);
        
    
        and(andpr47[10],b[46],a[10]);
        
    
        and(andpr47[11],b[46],a[11]);
        
    
        and(andpr47[12],b[46],a[12]);
        
    
        and(andpr47[13],b[46],a[13]);
        
    
        and(andpr47[14],b[46],a[14]);
        
    
        and(andpr47[15],b[46],a[15]);
        
    
        and(andpr47[16],b[46],a[16]);
        
    
        and(andpr47[17],b[46],a[17]);
        
    
        and(andpr47[18],b[46],a[18]);
        
    
        and(andpr47[19],b[46],a[19]);
        
    
        and(andpr47[20],b[46],a[20]);
        
    
        and(andpr47[21],b[46],a[21]);
        
    
        and(andpr47[22],b[46],a[22]);
        
    
        and(andpr47[23],b[46],a[23]);
        
    
        and(andpr47[24],b[46],a[24]);
        
    
        and(andpr47[25],b[46],a[25]);
        
    
        and(andpr47[26],b[46],a[26]);
        
    
        and(andpr47[27],b[46],a[27]);
        
    
        and(andpr47[28],b[46],a[28]);
        
    
        and(andpr47[29],b[46],a[29]);
        
    
        and(andpr47[30],b[46],a[30]);
        
    
        and(andpr47[31],b[46],a[31]);
        
    
        and(andpr47[32],b[46],a[32]);
        
    
        and(andpr47[33],b[46],a[33]);
        
    
        and(andpr47[34],b[46],a[34]);
        
    
        and(andpr47[35],b[46],a[35]);
        
    
        and(andpr47[36],b[46],a[36]);
        
    
        and(andpr47[37],b[46],a[37]);
        
    
        and(andpr47[38],b[46],a[38]);
        
    
        and(andpr47[39],b[46],a[39]);
        
    
        and(andpr47[40],b[46],a[40]);
        
    
        and(andpr47[41],b[46],a[41]);
        
    
        and(andpr47[42],b[46],a[42]);
        
    
        and(andpr47[43],b[46],a[43]);
        
    
        and(andpr47[44],b[46],a[44]);
        
    
        and(andpr47[45],b[46],a[45]);
        
    
        and(andpr47[46],b[46],a[46]);
        
    
        and(andpr47[47],b[46],a[47]);
        
    
        and(andpr47[48],b[46],a[48]);
        
    
        and(andpr47[49],b[46],a[49]);
        
    
        and(andpr47[50],b[46],a[50]);
        
    
        and(andpr47[51],b[46],a[51]);
        
    
        and(andpr47[52],b[46],a[52]);
        
    
        and(andpr47[53],b[46],a[53]);
        
    
        and(andpr47[54],b[46],a[54]);
        
    
        and(andpr47[55],b[46],a[55]);
        
    
        and(andpr47[56],b[46],a[56]);
        
    
        and(andpr47[57],b[46],a[57]);
        
    
        and(andpr47[58],b[46],a[58]);
        
    
        and(andpr47[59],b[46],a[59]);
        
    
        and(andpr47[60],b[46],a[60]);
        
    
        and(andpr47[61],b[46],a[61]);
        
    
        and(andpr47[62],b[46],a[62]);
        
    
        and(andpr47[63],b[46],a[63]);
        
    
    not(si[46],andpr47[63]);

    
        and(andpr48[0],b[47],a[0]);
        
    
        and(andpr48[1],b[47],a[1]);
        
    
        and(andpr48[2],b[47],a[2]);
        
    
        and(andpr48[3],b[47],a[3]);
        
    
        and(andpr48[4],b[47],a[4]);
        
    
        and(andpr48[5],b[47],a[5]);
        
    
        and(andpr48[6],b[47],a[6]);
        
    
        and(andpr48[7],b[47],a[7]);
        
    
        and(andpr48[8],b[47],a[8]);
        
    
        and(andpr48[9],b[47],a[9]);
        
    
        and(andpr48[10],b[47],a[10]);
        
    
        and(andpr48[11],b[47],a[11]);
        
    
        and(andpr48[12],b[47],a[12]);
        
    
        and(andpr48[13],b[47],a[13]);
        
    
        and(andpr48[14],b[47],a[14]);
        
    
        and(andpr48[15],b[47],a[15]);
        
    
        and(andpr48[16],b[47],a[16]);
        
    
        and(andpr48[17],b[47],a[17]);
        
    
        and(andpr48[18],b[47],a[18]);
        
    
        and(andpr48[19],b[47],a[19]);
        
    
        and(andpr48[20],b[47],a[20]);
        
    
        and(andpr48[21],b[47],a[21]);
        
    
        and(andpr48[22],b[47],a[22]);
        
    
        and(andpr48[23],b[47],a[23]);
        
    
        and(andpr48[24],b[47],a[24]);
        
    
        and(andpr48[25],b[47],a[25]);
        
    
        and(andpr48[26],b[47],a[26]);
        
    
        and(andpr48[27],b[47],a[27]);
        
    
        and(andpr48[28],b[47],a[28]);
        
    
        and(andpr48[29],b[47],a[29]);
        
    
        and(andpr48[30],b[47],a[30]);
        
    
        and(andpr48[31],b[47],a[31]);
        
    
        and(andpr48[32],b[47],a[32]);
        
    
        and(andpr48[33],b[47],a[33]);
        
    
        and(andpr48[34],b[47],a[34]);
        
    
        and(andpr48[35],b[47],a[35]);
        
    
        and(andpr48[36],b[47],a[36]);
        
    
        and(andpr48[37],b[47],a[37]);
        
    
        and(andpr48[38],b[47],a[38]);
        
    
        and(andpr48[39],b[47],a[39]);
        
    
        and(andpr48[40],b[47],a[40]);
        
    
        and(andpr48[41],b[47],a[41]);
        
    
        and(andpr48[42],b[47],a[42]);
        
    
        and(andpr48[43],b[47],a[43]);
        
    
        and(andpr48[44],b[47],a[44]);
        
    
        and(andpr48[45],b[47],a[45]);
        
    
        and(andpr48[46],b[47],a[46]);
        
    
        and(andpr48[47],b[47],a[47]);
        
    
        and(andpr48[48],b[47],a[48]);
        
    
        and(andpr48[49],b[47],a[49]);
        
    
        and(andpr48[50],b[47],a[50]);
        
    
        and(andpr48[51],b[47],a[51]);
        
    
        and(andpr48[52],b[47],a[52]);
        
    
        and(andpr48[53],b[47],a[53]);
        
    
        and(andpr48[54],b[47],a[54]);
        
    
        and(andpr48[55],b[47],a[55]);
        
    
        and(andpr48[56],b[47],a[56]);
        
    
        and(andpr48[57],b[47],a[57]);
        
    
        and(andpr48[58],b[47],a[58]);
        
    
        and(andpr48[59],b[47],a[59]);
        
    
        and(andpr48[60],b[47],a[60]);
        
    
        and(andpr48[61],b[47],a[61]);
        
    
        and(andpr48[62],b[47],a[62]);
        
    
        and(andpr48[63],b[47],a[63]);
        
    
    not(si[47],andpr48[63]);

    
        and(andpr49[0],b[48],a[0]);
        
    
        and(andpr49[1],b[48],a[1]);
        
    
        and(andpr49[2],b[48],a[2]);
        
    
        and(andpr49[3],b[48],a[3]);
        
    
        and(andpr49[4],b[48],a[4]);
        
    
        and(andpr49[5],b[48],a[5]);
        
    
        and(andpr49[6],b[48],a[6]);
        
    
        and(andpr49[7],b[48],a[7]);
        
    
        and(andpr49[8],b[48],a[8]);
        
    
        and(andpr49[9],b[48],a[9]);
        
    
        and(andpr49[10],b[48],a[10]);
        
    
        and(andpr49[11],b[48],a[11]);
        
    
        and(andpr49[12],b[48],a[12]);
        
    
        and(andpr49[13],b[48],a[13]);
        
    
        and(andpr49[14],b[48],a[14]);
        
    
        and(andpr49[15],b[48],a[15]);
        
    
        and(andpr49[16],b[48],a[16]);
        
    
        and(andpr49[17],b[48],a[17]);
        
    
        and(andpr49[18],b[48],a[18]);
        
    
        and(andpr49[19],b[48],a[19]);
        
    
        and(andpr49[20],b[48],a[20]);
        
    
        and(andpr49[21],b[48],a[21]);
        
    
        and(andpr49[22],b[48],a[22]);
        
    
        and(andpr49[23],b[48],a[23]);
        
    
        and(andpr49[24],b[48],a[24]);
        
    
        and(andpr49[25],b[48],a[25]);
        
    
        and(andpr49[26],b[48],a[26]);
        
    
        and(andpr49[27],b[48],a[27]);
        
    
        and(andpr49[28],b[48],a[28]);
        
    
        and(andpr49[29],b[48],a[29]);
        
    
        and(andpr49[30],b[48],a[30]);
        
    
        and(andpr49[31],b[48],a[31]);
        
    
        and(andpr49[32],b[48],a[32]);
        
    
        and(andpr49[33],b[48],a[33]);
        
    
        and(andpr49[34],b[48],a[34]);
        
    
        and(andpr49[35],b[48],a[35]);
        
    
        and(andpr49[36],b[48],a[36]);
        
    
        and(andpr49[37],b[48],a[37]);
        
    
        and(andpr49[38],b[48],a[38]);
        
    
        and(andpr49[39],b[48],a[39]);
        
    
        and(andpr49[40],b[48],a[40]);
        
    
        and(andpr49[41],b[48],a[41]);
        
    
        and(andpr49[42],b[48],a[42]);
        
    
        and(andpr49[43],b[48],a[43]);
        
    
        and(andpr49[44],b[48],a[44]);
        
    
        and(andpr49[45],b[48],a[45]);
        
    
        and(andpr49[46],b[48],a[46]);
        
    
        and(andpr49[47],b[48],a[47]);
        
    
        and(andpr49[48],b[48],a[48]);
        
    
        and(andpr49[49],b[48],a[49]);
        
    
        and(andpr49[50],b[48],a[50]);
        
    
        and(andpr49[51],b[48],a[51]);
        
    
        and(andpr49[52],b[48],a[52]);
        
    
        and(andpr49[53],b[48],a[53]);
        
    
        and(andpr49[54],b[48],a[54]);
        
    
        and(andpr49[55],b[48],a[55]);
        
    
        and(andpr49[56],b[48],a[56]);
        
    
        and(andpr49[57],b[48],a[57]);
        
    
        and(andpr49[58],b[48],a[58]);
        
    
        and(andpr49[59],b[48],a[59]);
        
    
        and(andpr49[60],b[48],a[60]);
        
    
        and(andpr49[61],b[48],a[61]);
        
    
        and(andpr49[62],b[48],a[62]);
        
    
        and(andpr49[63],b[48],a[63]);
        
    
    not(si[48],andpr49[63]);

    
        and(andpr50[0],b[49],a[0]);
        
    
        and(andpr50[1],b[49],a[1]);
        
    
        and(andpr50[2],b[49],a[2]);
        
    
        and(andpr50[3],b[49],a[3]);
        
    
        and(andpr50[4],b[49],a[4]);
        
    
        and(andpr50[5],b[49],a[5]);
        
    
        and(andpr50[6],b[49],a[6]);
        
    
        and(andpr50[7],b[49],a[7]);
        
    
        and(andpr50[8],b[49],a[8]);
        
    
        and(andpr50[9],b[49],a[9]);
        
    
        and(andpr50[10],b[49],a[10]);
        
    
        and(andpr50[11],b[49],a[11]);
        
    
        and(andpr50[12],b[49],a[12]);
        
    
        and(andpr50[13],b[49],a[13]);
        
    
        and(andpr50[14],b[49],a[14]);
        
    
        and(andpr50[15],b[49],a[15]);
        
    
        and(andpr50[16],b[49],a[16]);
        
    
        and(andpr50[17],b[49],a[17]);
        
    
        and(andpr50[18],b[49],a[18]);
        
    
        and(andpr50[19],b[49],a[19]);
        
    
        and(andpr50[20],b[49],a[20]);
        
    
        and(andpr50[21],b[49],a[21]);
        
    
        and(andpr50[22],b[49],a[22]);
        
    
        and(andpr50[23],b[49],a[23]);
        
    
        and(andpr50[24],b[49],a[24]);
        
    
        and(andpr50[25],b[49],a[25]);
        
    
        and(andpr50[26],b[49],a[26]);
        
    
        and(andpr50[27],b[49],a[27]);
        
    
        and(andpr50[28],b[49],a[28]);
        
    
        and(andpr50[29],b[49],a[29]);
        
    
        and(andpr50[30],b[49],a[30]);
        
    
        and(andpr50[31],b[49],a[31]);
        
    
        and(andpr50[32],b[49],a[32]);
        
    
        and(andpr50[33],b[49],a[33]);
        
    
        and(andpr50[34],b[49],a[34]);
        
    
        and(andpr50[35],b[49],a[35]);
        
    
        and(andpr50[36],b[49],a[36]);
        
    
        and(andpr50[37],b[49],a[37]);
        
    
        and(andpr50[38],b[49],a[38]);
        
    
        and(andpr50[39],b[49],a[39]);
        
    
        and(andpr50[40],b[49],a[40]);
        
    
        and(andpr50[41],b[49],a[41]);
        
    
        and(andpr50[42],b[49],a[42]);
        
    
        and(andpr50[43],b[49],a[43]);
        
    
        and(andpr50[44],b[49],a[44]);
        
    
        and(andpr50[45],b[49],a[45]);
        
    
        and(andpr50[46],b[49],a[46]);
        
    
        and(andpr50[47],b[49],a[47]);
        
    
        and(andpr50[48],b[49],a[48]);
        
    
        and(andpr50[49],b[49],a[49]);
        
    
        and(andpr50[50],b[49],a[50]);
        
    
        and(andpr50[51],b[49],a[51]);
        
    
        and(andpr50[52],b[49],a[52]);
        
    
        and(andpr50[53],b[49],a[53]);
        
    
        and(andpr50[54],b[49],a[54]);
        
    
        and(andpr50[55],b[49],a[55]);
        
    
        and(andpr50[56],b[49],a[56]);
        
    
        and(andpr50[57],b[49],a[57]);
        
    
        and(andpr50[58],b[49],a[58]);
        
    
        and(andpr50[59],b[49],a[59]);
        
    
        and(andpr50[60],b[49],a[60]);
        
    
        and(andpr50[61],b[49],a[61]);
        
    
        and(andpr50[62],b[49],a[62]);
        
    
        and(andpr50[63],b[49],a[63]);
        
    
    not(si[49],andpr50[63]);

    
        and(andpr51[0],b[50],a[0]);
        
    
        and(andpr51[1],b[50],a[1]);
        
    
        and(andpr51[2],b[50],a[2]);
        
    
        and(andpr51[3],b[50],a[3]);
        
    
        and(andpr51[4],b[50],a[4]);
        
    
        and(andpr51[5],b[50],a[5]);
        
    
        and(andpr51[6],b[50],a[6]);
        
    
        and(andpr51[7],b[50],a[7]);
        
    
        and(andpr51[8],b[50],a[8]);
        
    
        and(andpr51[9],b[50],a[9]);
        
    
        and(andpr51[10],b[50],a[10]);
        
    
        and(andpr51[11],b[50],a[11]);
        
    
        and(andpr51[12],b[50],a[12]);
        
    
        and(andpr51[13],b[50],a[13]);
        
    
        and(andpr51[14],b[50],a[14]);
        
    
        and(andpr51[15],b[50],a[15]);
        
    
        and(andpr51[16],b[50],a[16]);
        
    
        and(andpr51[17],b[50],a[17]);
        
    
        and(andpr51[18],b[50],a[18]);
        
    
        and(andpr51[19],b[50],a[19]);
        
    
        and(andpr51[20],b[50],a[20]);
        
    
        and(andpr51[21],b[50],a[21]);
        
    
        and(andpr51[22],b[50],a[22]);
        
    
        and(andpr51[23],b[50],a[23]);
        
    
        and(andpr51[24],b[50],a[24]);
        
    
        and(andpr51[25],b[50],a[25]);
        
    
        and(andpr51[26],b[50],a[26]);
        
    
        and(andpr51[27],b[50],a[27]);
        
    
        and(andpr51[28],b[50],a[28]);
        
    
        and(andpr51[29],b[50],a[29]);
        
    
        and(andpr51[30],b[50],a[30]);
        
    
        and(andpr51[31],b[50],a[31]);
        
    
        and(andpr51[32],b[50],a[32]);
        
    
        and(andpr51[33],b[50],a[33]);
        
    
        and(andpr51[34],b[50],a[34]);
        
    
        and(andpr51[35],b[50],a[35]);
        
    
        and(andpr51[36],b[50],a[36]);
        
    
        and(andpr51[37],b[50],a[37]);
        
    
        and(andpr51[38],b[50],a[38]);
        
    
        and(andpr51[39],b[50],a[39]);
        
    
        and(andpr51[40],b[50],a[40]);
        
    
        and(andpr51[41],b[50],a[41]);
        
    
        and(andpr51[42],b[50],a[42]);
        
    
        and(andpr51[43],b[50],a[43]);
        
    
        and(andpr51[44],b[50],a[44]);
        
    
        and(andpr51[45],b[50],a[45]);
        
    
        and(andpr51[46],b[50],a[46]);
        
    
        and(andpr51[47],b[50],a[47]);
        
    
        and(andpr51[48],b[50],a[48]);
        
    
        and(andpr51[49],b[50],a[49]);
        
    
        and(andpr51[50],b[50],a[50]);
        
    
        and(andpr51[51],b[50],a[51]);
        
    
        and(andpr51[52],b[50],a[52]);
        
    
        and(andpr51[53],b[50],a[53]);
        
    
        and(andpr51[54],b[50],a[54]);
        
    
        and(andpr51[55],b[50],a[55]);
        
    
        and(andpr51[56],b[50],a[56]);
        
    
        and(andpr51[57],b[50],a[57]);
        
    
        and(andpr51[58],b[50],a[58]);
        
    
        and(andpr51[59],b[50],a[59]);
        
    
        and(andpr51[60],b[50],a[60]);
        
    
        and(andpr51[61],b[50],a[61]);
        
    
        and(andpr51[62],b[50],a[62]);
        
    
        and(andpr51[63],b[50],a[63]);
        
    
    not(si[50],andpr51[63]);

    
        and(andpr52[0],b[51],a[0]);
        
    
        and(andpr52[1],b[51],a[1]);
        
    
        and(andpr52[2],b[51],a[2]);
        
    
        and(andpr52[3],b[51],a[3]);
        
    
        and(andpr52[4],b[51],a[4]);
        
    
        and(andpr52[5],b[51],a[5]);
        
    
        and(andpr52[6],b[51],a[6]);
        
    
        and(andpr52[7],b[51],a[7]);
        
    
        and(andpr52[8],b[51],a[8]);
        
    
        and(andpr52[9],b[51],a[9]);
        
    
        and(andpr52[10],b[51],a[10]);
        
    
        and(andpr52[11],b[51],a[11]);
        
    
        and(andpr52[12],b[51],a[12]);
        
    
        and(andpr52[13],b[51],a[13]);
        
    
        and(andpr52[14],b[51],a[14]);
        
    
        and(andpr52[15],b[51],a[15]);
        
    
        and(andpr52[16],b[51],a[16]);
        
    
        and(andpr52[17],b[51],a[17]);
        
    
        and(andpr52[18],b[51],a[18]);
        
    
        and(andpr52[19],b[51],a[19]);
        
    
        and(andpr52[20],b[51],a[20]);
        
    
        and(andpr52[21],b[51],a[21]);
        
    
        and(andpr52[22],b[51],a[22]);
        
    
        and(andpr52[23],b[51],a[23]);
        
    
        and(andpr52[24],b[51],a[24]);
        
    
        and(andpr52[25],b[51],a[25]);
        
    
        and(andpr52[26],b[51],a[26]);
        
    
        and(andpr52[27],b[51],a[27]);
        
    
        and(andpr52[28],b[51],a[28]);
        
    
        and(andpr52[29],b[51],a[29]);
        
    
        and(andpr52[30],b[51],a[30]);
        
    
        and(andpr52[31],b[51],a[31]);
        
    
        and(andpr52[32],b[51],a[32]);
        
    
        and(andpr52[33],b[51],a[33]);
        
    
        and(andpr52[34],b[51],a[34]);
        
    
        and(andpr52[35],b[51],a[35]);
        
    
        and(andpr52[36],b[51],a[36]);
        
    
        and(andpr52[37],b[51],a[37]);
        
    
        and(andpr52[38],b[51],a[38]);
        
    
        and(andpr52[39],b[51],a[39]);
        
    
        and(andpr52[40],b[51],a[40]);
        
    
        and(andpr52[41],b[51],a[41]);
        
    
        and(andpr52[42],b[51],a[42]);
        
    
        and(andpr52[43],b[51],a[43]);
        
    
        and(andpr52[44],b[51],a[44]);
        
    
        and(andpr52[45],b[51],a[45]);
        
    
        and(andpr52[46],b[51],a[46]);
        
    
        and(andpr52[47],b[51],a[47]);
        
    
        and(andpr52[48],b[51],a[48]);
        
    
        and(andpr52[49],b[51],a[49]);
        
    
        and(andpr52[50],b[51],a[50]);
        
    
        and(andpr52[51],b[51],a[51]);
        
    
        and(andpr52[52],b[51],a[52]);
        
    
        and(andpr52[53],b[51],a[53]);
        
    
        and(andpr52[54],b[51],a[54]);
        
    
        and(andpr52[55],b[51],a[55]);
        
    
        and(andpr52[56],b[51],a[56]);
        
    
        and(andpr52[57],b[51],a[57]);
        
    
        and(andpr52[58],b[51],a[58]);
        
    
        and(andpr52[59],b[51],a[59]);
        
    
        and(andpr52[60],b[51],a[60]);
        
    
        and(andpr52[61],b[51],a[61]);
        
    
        and(andpr52[62],b[51],a[62]);
        
    
        and(andpr52[63],b[51],a[63]);
        
    
    not(si[51],andpr52[63]);

    
        and(andpr53[0],b[52],a[0]);
        
    
        and(andpr53[1],b[52],a[1]);
        
    
        and(andpr53[2],b[52],a[2]);
        
    
        and(andpr53[3],b[52],a[3]);
        
    
        and(andpr53[4],b[52],a[4]);
        
    
        and(andpr53[5],b[52],a[5]);
        
    
        and(andpr53[6],b[52],a[6]);
        
    
        and(andpr53[7],b[52],a[7]);
        
    
        and(andpr53[8],b[52],a[8]);
        
    
        and(andpr53[9],b[52],a[9]);
        
    
        and(andpr53[10],b[52],a[10]);
        
    
        and(andpr53[11],b[52],a[11]);
        
    
        and(andpr53[12],b[52],a[12]);
        
    
        and(andpr53[13],b[52],a[13]);
        
    
        and(andpr53[14],b[52],a[14]);
        
    
        and(andpr53[15],b[52],a[15]);
        
    
        and(andpr53[16],b[52],a[16]);
        
    
        and(andpr53[17],b[52],a[17]);
        
    
        and(andpr53[18],b[52],a[18]);
        
    
        and(andpr53[19],b[52],a[19]);
        
    
        and(andpr53[20],b[52],a[20]);
        
    
        and(andpr53[21],b[52],a[21]);
        
    
        and(andpr53[22],b[52],a[22]);
        
    
        and(andpr53[23],b[52],a[23]);
        
    
        and(andpr53[24],b[52],a[24]);
        
    
        and(andpr53[25],b[52],a[25]);
        
    
        and(andpr53[26],b[52],a[26]);
        
    
        and(andpr53[27],b[52],a[27]);
        
    
        and(andpr53[28],b[52],a[28]);
        
    
        and(andpr53[29],b[52],a[29]);
        
    
        and(andpr53[30],b[52],a[30]);
        
    
        and(andpr53[31],b[52],a[31]);
        
    
        and(andpr53[32],b[52],a[32]);
        
    
        and(andpr53[33],b[52],a[33]);
        
    
        and(andpr53[34],b[52],a[34]);
        
    
        and(andpr53[35],b[52],a[35]);
        
    
        and(andpr53[36],b[52],a[36]);
        
    
        and(andpr53[37],b[52],a[37]);
        
    
        and(andpr53[38],b[52],a[38]);
        
    
        and(andpr53[39],b[52],a[39]);
        
    
        and(andpr53[40],b[52],a[40]);
        
    
        and(andpr53[41],b[52],a[41]);
        
    
        and(andpr53[42],b[52],a[42]);
        
    
        and(andpr53[43],b[52],a[43]);
        
    
        and(andpr53[44],b[52],a[44]);
        
    
        and(andpr53[45],b[52],a[45]);
        
    
        and(andpr53[46],b[52],a[46]);
        
    
        and(andpr53[47],b[52],a[47]);
        
    
        and(andpr53[48],b[52],a[48]);
        
    
        and(andpr53[49],b[52],a[49]);
        
    
        and(andpr53[50],b[52],a[50]);
        
    
        and(andpr53[51],b[52],a[51]);
        
    
        and(andpr53[52],b[52],a[52]);
        
    
        and(andpr53[53],b[52],a[53]);
        
    
        and(andpr53[54],b[52],a[54]);
        
    
        and(andpr53[55],b[52],a[55]);
        
    
        and(andpr53[56],b[52],a[56]);
        
    
        and(andpr53[57],b[52],a[57]);
        
    
        and(andpr53[58],b[52],a[58]);
        
    
        and(andpr53[59],b[52],a[59]);
        
    
        and(andpr53[60],b[52],a[60]);
        
    
        and(andpr53[61],b[52],a[61]);
        
    
        and(andpr53[62],b[52],a[62]);
        
    
        and(andpr53[63],b[52],a[63]);
        
    
    not(si[52],andpr53[63]);

    
        and(andpr54[0],b[53],a[0]);
        
    
        and(andpr54[1],b[53],a[1]);
        
    
        and(andpr54[2],b[53],a[2]);
        
    
        and(andpr54[3],b[53],a[3]);
        
    
        and(andpr54[4],b[53],a[4]);
        
    
        and(andpr54[5],b[53],a[5]);
        
    
        and(andpr54[6],b[53],a[6]);
        
    
        and(andpr54[7],b[53],a[7]);
        
    
        and(andpr54[8],b[53],a[8]);
        
    
        and(andpr54[9],b[53],a[9]);
        
    
        and(andpr54[10],b[53],a[10]);
        
    
        and(andpr54[11],b[53],a[11]);
        
    
        and(andpr54[12],b[53],a[12]);
        
    
        and(andpr54[13],b[53],a[13]);
        
    
        and(andpr54[14],b[53],a[14]);
        
    
        and(andpr54[15],b[53],a[15]);
        
    
        and(andpr54[16],b[53],a[16]);
        
    
        and(andpr54[17],b[53],a[17]);
        
    
        and(andpr54[18],b[53],a[18]);
        
    
        and(andpr54[19],b[53],a[19]);
        
    
        and(andpr54[20],b[53],a[20]);
        
    
        and(andpr54[21],b[53],a[21]);
        
    
        and(andpr54[22],b[53],a[22]);
        
    
        and(andpr54[23],b[53],a[23]);
        
    
        and(andpr54[24],b[53],a[24]);
        
    
        and(andpr54[25],b[53],a[25]);
        
    
        and(andpr54[26],b[53],a[26]);
        
    
        and(andpr54[27],b[53],a[27]);
        
    
        and(andpr54[28],b[53],a[28]);
        
    
        and(andpr54[29],b[53],a[29]);
        
    
        and(andpr54[30],b[53],a[30]);
        
    
        and(andpr54[31],b[53],a[31]);
        
    
        and(andpr54[32],b[53],a[32]);
        
    
        and(andpr54[33],b[53],a[33]);
        
    
        and(andpr54[34],b[53],a[34]);
        
    
        and(andpr54[35],b[53],a[35]);
        
    
        and(andpr54[36],b[53],a[36]);
        
    
        and(andpr54[37],b[53],a[37]);
        
    
        and(andpr54[38],b[53],a[38]);
        
    
        and(andpr54[39],b[53],a[39]);
        
    
        and(andpr54[40],b[53],a[40]);
        
    
        and(andpr54[41],b[53],a[41]);
        
    
        and(andpr54[42],b[53],a[42]);
        
    
        and(andpr54[43],b[53],a[43]);
        
    
        and(andpr54[44],b[53],a[44]);
        
    
        and(andpr54[45],b[53],a[45]);
        
    
        and(andpr54[46],b[53],a[46]);
        
    
        and(andpr54[47],b[53],a[47]);
        
    
        and(andpr54[48],b[53],a[48]);
        
    
        and(andpr54[49],b[53],a[49]);
        
    
        and(andpr54[50],b[53],a[50]);
        
    
        and(andpr54[51],b[53],a[51]);
        
    
        and(andpr54[52],b[53],a[52]);
        
    
        and(andpr54[53],b[53],a[53]);
        
    
        and(andpr54[54],b[53],a[54]);
        
    
        and(andpr54[55],b[53],a[55]);
        
    
        and(andpr54[56],b[53],a[56]);
        
    
        and(andpr54[57],b[53],a[57]);
        
    
        and(andpr54[58],b[53],a[58]);
        
    
        and(andpr54[59],b[53],a[59]);
        
    
        and(andpr54[60],b[53],a[60]);
        
    
        and(andpr54[61],b[53],a[61]);
        
    
        and(andpr54[62],b[53],a[62]);
        
    
        and(andpr54[63],b[53],a[63]);
        
    
    not(si[53],andpr54[63]);

    
        and(andpr55[0],b[54],a[0]);
        
    
        and(andpr55[1],b[54],a[1]);
        
    
        and(andpr55[2],b[54],a[2]);
        
    
        and(andpr55[3],b[54],a[3]);
        
    
        and(andpr55[4],b[54],a[4]);
        
    
        and(andpr55[5],b[54],a[5]);
        
    
        and(andpr55[6],b[54],a[6]);
        
    
        and(andpr55[7],b[54],a[7]);
        
    
        and(andpr55[8],b[54],a[8]);
        
    
        and(andpr55[9],b[54],a[9]);
        
    
        and(andpr55[10],b[54],a[10]);
        
    
        and(andpr55[11],b[54],a[11]);
        
    
        and(andpr55[12],b[54],a[12]);
        
    
        and(andpr55[13],b[54],a[13]);
        
    
        and(andpr55[14],b[54],a[14]);
        
    
        and(andpr55[15],b[54],a[15]);
        
    
        and(andpr55[16],b[54],a[16]);
        
    
        and(andpr55[17],b[54],a[17]);
        
    
        and(andpr55[18],b[54],a[18]);
        
    
        and(andpr55[19],b[54],a[19]);
        
    
        and(andpr55[20],b[54],a[20]);
        
    
        and(andpr55[21],b[54],a[21]);
        
    
        and(andpr55[22],b[54],a[22]);
        
    
        and(andpr55[23],b[54],a[23]);
        
    
        and(andpr55[24],b[54],a[24]);
        
    
        and(andpr55[25],b[54],a[25]);
        
    
        and(andpr55[26],b[54],a[26]);
        
    
        and(andpr55[27],b[54],a[27]);
        
    
        and(andpr55[28],b[54],a[28]);
        
    
        and(andpr55[29],b[54],a[29]);
        
    
        and(andpr55[30],b[54],a[30]);
        
    
        and(andpr55[31],b[54],a[31]);
        
    
        and(andpr55[32],b[54],a[32]);
        
    
        and(andpr55[33],b[54],a[33]);
        
    
        and(andpr55[34],b[54],a[34]);
        
    
        and(andpr55[35],b[54],a[35]);
        
    
        and(andpr55[36],b[54],a[36]);
        
    
        and(andpr55[37],b[54],a[37]);
        
    
        and(andpr55[38],b[54],a[38]);
        
    
        and(andpr55[39],b[54],a[39]);
        
    
        and(andpr55[40],b[54],a[40]);
        
    
        and(andpr55[41],b[54],a[41]);
        
    
        and(andpr55[42],b[54],a[42]);
        
    
        and(andpr55[43],b[54],a[43]);
        
    
        and(andpr55[44],b[54],a[44]);
        
    
        and(andpr55[45],b[54],a[45]);
        
    
        and(andpr55[46],b[54],a[46]);
        
    
        and(andpr55[47],b[54],a[47]);
        
    
        and(andpr55[48],b[54],a[48]);
        
    
        and(andpr55[49],b[54],a[49]);
        
    
        and(andpr55[50],b[54],a[50]);
        
    
        and(andpr55[51],b[54],a[51]);
        
    
        and(andpr55[52],b[54],a[52]);
        
    
        and(andpr55[53],b[54],a[53]);
        
    
        and(andpr55[54],b[54],a[54]);
        
    
        and(andpr55[55],b[54],a[55]);
        
    
        and(andpr55[56],b[54],a[56]);
        
    
        and(andpr55[57],b[54],a[57]);
        
    
        and(andpr55[58],b[54],a[58]);
        
    
        and(andpr55[59],b[54],a[59]);
        
    
        and(andpr55[60],b[54],a[60]);
        
    
        and(andpr55[61],b[54],a[61]);
        
    
        and(andpr55[62],b[54],a[62]);
        
    
        and(andpr55[63],b[54],a[63]);
        
    
    not(si[54],andpr55[63]);

    
        and(andpr56[0],b[55],a[0]);
        
    
        and(andpr56[1],b[55],a[1]);
        
    
        and(andpr56[2],b[55],a[2]);
        
    
        and(andpr56[3],b[55],a[3]);
        
    
        and(andpr56[4],b[55],a[4]);
        
    
        and(andpr56[5],b[55],a[5]);
        
    
        and(andpr56[6],b[55],a[6]);
        
    
        and(andpr56[7],b[55],a[7]);
        
    
        and(andpr56[8],b[55],a[8]);
        
    
        and(andpr56[9],b[55],a[9]);
        
    
        and(andpr56[10],b[55],a[10]);
        
    
        and(andpr56[11],b[55],a[11]);
        
    
        and(andpr56[12],b[55],a[12]);
        
    
        and(andpr56[13],b[55],a[13]);
        
    
        and(andpr56[14],b[55],a[14]);
        
    
        and(andpr56[15],b[55],a[15]);
        
    
        and(andpr56[16],b[55],a[16]);
        
    
        and(andpr56[17],b[55],a[17]);
        
    
        and(andpr56[18],b[55],a[18]);
        
    
        and(andpr56[19],b[55],a[19]);
        
    
        and(andpr56[20],b[55],a[20]);
        
    
        and(andpr56[21],b[55],a[21]);
        
    
        and(andpr56[22],b[55],a[22]);
        
    
        and(andpr56[23],b[55],a[23]);
        
    
        and(andpr56[24],b[55],a[24]);
        
    
        and(andpr56[25],b[55],a[25]);
        
    
        and(andpr56[26],b[55],a[26]);
        
    
        and(andpr56[27],b[55],a[27]);
        
    
        and(andpr56[28],b[55],a[28]);
        
    
        and(andpr56[29],b[55],a[29]);
        
    
        and(andpr56[30],b[55],a[30]);
        
    
        and(andpr56[31],b[55],a[31]);
        
    
        and(andpr56[32],b[55],a[32]);
        
    
        and(andpr56[33],b[55],a[33]);
        
    
        and(andpr56[34],b[55],a[34]);
        
    
        and(andpr56[35],b[55],a[35]);
        
    
        and(andpr56[36],b[55],a[36]);
        
    
        and(andpr56[37],b[55],a[37]);
        
    
        and(andpr56[38],b[55],a[38]);
        
    
        and(andpr56[39],b[55],a[39]);
        
    
        and(andpr56[40],b[55],a[40]);
        
    
        and(andpr56[41],b[55],a[41]);
        
    
        and(andpr56[42],b[55],a[42]);
        
    
        and(andpr56[43],b[55],a[43]);
        
    
        and(andpr56[44],b[55],a[44]);
        
    
        and(andpr56[45],b[55],a[45]);
        
    
        and(andpr56[46],b[55],a[46]);
        
    
        and(andpr56[47],b[55],a[47]);
        
    
        and(andpr56[48],b[55],a[48]);
        
    
        and(andpr56[49],b[55],a[49]);
        
    
        and(andpr56[50],b[55],a[50]);
        
    
        and(andpr56[51],b[55],a[51]);
        
    
        and(andpr56[52],b[55],a[52]);
        
    
        and(andpr56[53],b[55],a[53]);
        
    
        and(andpr56[54],b[55],a[54]);
        
    
        and(andpr56[55],b[55],a[55]);
        
    
        and(andpr56[56],b[55],a[56]);
        
    
        and(andpr56[57],b[55],a[57]);
        
    
        and(andpr56[58],b[55],a[58]);
        
    
        and(andpr56[59],b[55],a[59]);
        
    
        and(andpr56[60],b[55],a[60]);
        
    
        and(andpr56[61],b[55],a[61]);
        
    
        and(andpr56[62],b[55],a[62]);
        
    
        and(andpr56[63],b[55],a[63]);
        
    
    not(si[55],andpr56[63]);

    
        and(andpr57[0],b[56],a[0]);
        
    
        and(andpr57[1],b[56],a[1]);
        
    
        and(andpr57[2],b[56],a[2]);
        
    
        and(andpr57[3],b[56],a[3]);
        
    
        and(andpr57[4],b[56],a[4]);
        
    
        and(andpr57[5],b[56],a[5]);
        
    
        and(andpr57[6],b[56],a[6]);
        
    
        and(andpr57[7],b[56],a[7]);
        
    
        and(andpr57[8],b[56],a[8]);
        
    
        and(andpr57[9],b[56],a[9]);
        
    
        and(andpr57[10],b[56],a[10]);
        
    
        and(andpr57[11],b[56],a[11]);
        
    
        and(andpr57[12],b[56],a[12]);
        
    
        and(andpr57[13],b[56],a[13]);
        
    
        and(andpr57[14],b[56],a[14]);
        
    
        and(andpr57[15],b[56],a[15]);
        
    
        and(andpr57[16],b[56],a[16]);
        
    
        and(andpr57[17],b[56],a[17]);
        
    
        and(andpr57[18],b[56],a[18]);
        
    
        and(andpr57[19],b[56],a[19]);
        
    
        and(andpr57[20],b[56],a[20]);
        
    
        and(andpr57[21],b[56],a[21]);
        
    
        and(andpr57[22],b[56],a[22]);
        
    
        and(andpr57[23],b[56],a[23]);
        
    
        and(andpr57[24],b[56],a[24]);
        
    
        and(andpr57[25],b[56],a[25]);
        
    
        and(andpr57[26],b[56],a[26]);
        
    
        and(andpr57[27],b[56],a[27]);
        
    
        and(andpr57[28],b[56],a[28]);
        
    
        and(andpr57[29],b[56],a[29]);
        
    
        and(andpr57[30],b[56],a[30]);
        
    
        and(andpr57[31],b[56],a[31]);
        
    
        and(andpr57[32],b[56],a[32]);
        
    
        and(andpr57[33],b[56],a[33]);
        
    
        and(andpr57[34],b[56],a[34]);
        
    
        and(andpr57[35],b[56],a[35]);
        
    
        and(andpr57[36],b[56],a[36]);
        
    
        and(andpr57[37],b[56],a[37]);
        
    
        and(andpr57[38],b[56],a[38]);
        
    
        and(andpr57[39],b[56],a[39]);
        
    
        and(andpr57[40],b[56],a[40]);
        
    
        and(andpr57[41],b[56],a[41]);
        
    
        and(andpr57[42],b[56],a[42]);
        
    
        and(andpr57[43],b[56],a[43]);
        
    
        and(andpr57[44],b[56],a[44]);
        
    
        and(andpr57[45],b[56],a[45]);
        
    
        and(andpr57[46],b[56],a[46]);
        
    
        and(andpr57[47],b[56],a[47]);
        
    
        and(andpr57[48],b[56],a[48]);
        
    
        and(andpr57[49],b[56],a[49]);
        
    
        and(andpr57[50],b[56],a[50]);
        
    
        and(andpr57[51],b[56],a[51]);
        
    
        and(andpr57[52],b[56],a[52]);
        
    
        and(andpr57[53],b[56],a[53]);
        
    
        and(andpr57[54],b[56],a[54]);
        
    
        and(andpr57[55],b[56],a[55]);
        
    
        and(andpr57[56],b[56],a[56]);
        
    
        and(andpr57[57],b[56],a[57]);
        
    
        and(andpr57[58],b[56],a[58]);
        
    
        and(andpr57[59],b[56],a[59]);
        
    
        and(andpr57[60],b[56],a[60]);
        
    
        and(andpr57[61],b[56],a[61]);
        
    
        and(andpr57[62],b[56],a[62]);
        
    
        and(andpr57[63],b[56],a[63]);
        
    
    not(si[56],andpr57[63]);

    
        and(andpr58[0],b[57],a[0]);
        
    
        and(andpr58[1],b[57],a[1]);
        
    
        and(andpr58[2],b[57],a[2]);
        
    
        and(andpr58[3],b[57],a[3]);
        
    
        and(andpr58[4],b[57],a[4]);
        
    
        and(andpr58[5],b[57],a[5]);
        
    
        and(andpr58[6],b[57],a[6]);
        
    
        and(andpr58[7],b[57],a[7]);
        
    
        and(andpr58[8],b[57],a[8]);
        
    
        and(andpr58[9],b[57],a[9]);
        
    
        and(andpr58[10],b[57],a[10]);
        
    
        and(andpr58[11],b[57],a[11]);
        
    
        and(andpr58[12],b[57],a[12]);
        
    
        and(andpr58[13],b[57],a[13]);
        
    
        and(andpr58[14],b[57],a[14]);
        
    
        and(andpr58[15],b[57],a[15]);
        
    
        and(andpr58[16],b[57],a[16]);
        
    
        and(andpr58[17],b[57],a[17]);
        
    
        and(andpr58[18],b[57],a[18]);
        
    
        and(andpr58[19],b[57],a[19]);
        
    
        and(andpr58[20],b[57],a[20]);
        
    
        and(andpr58[21],b[57],a[21]);
        
    
        and(andpr58[22],b[57],a[22]);
        
    
        and(andpr58[23],b[57],a[23]);
        
    
        and(andpr58[24],b[57],a[24]);
        
    
        and(andpr58[25],b[57],a[25]);
        
    
        and(andpr58[26],b[57],a[26]);
        
    
        and(andpr58[27],b[57],a[27]);
        
    
        and(andpr58[28],b[57],a[28]);
        
    
        and(andpr58[29],b[57],a[29]);
        
    
        and(andpr58[30],b[57],a[30]);
        
    
        and(andpr58[31],b[57],a[31]);
        
    
        and(andpr58[32],b[57],a[32]);
        
    
        and(andpr58[33],b[57],a[33]);
        
    
        and(andpr58[34],b[57],a[34]);
        
    
        and(andpr58[35],b[57],a[35]);
        
    
        and(andpr58[36],b[57],a[36]);
        
    
        and(andpr58[37],b[57],a[37]);
        
    
        and(andpr58[38],b[57],a[38]);
        
    
        and(andpr58[39],b[57],a[39]);
        
    
        and(andpr58[40],b[57],a[40]);
        
    
        and(andpr58[41],b[57],a[41]);
        
    
        and(andpr58[42],b[57],a[42]);
        
    
        and(andpr58[43],b[57],a[43]);
        
    
        and(andpr58[44],b[57],a[44]);
        
    
        and(andpr58[45],b[57],a[45]);
        
    
        and(andpr58[46],b[57],a[46]);
        
    
        and(andpr58[47],b[57],a[47]);
        
    
        and(andpr58[48],b[57],a[48]);
        
    
        and(andpr58[49],b[57],a[49]);
        
    
        and(andpr58[50],b[57],a[50]);
        
    
        and(andpr58[51],b[57],a[51]);
        
    
        and(andpr58[52],b[57],a[52]);
        
    
        and(andpr58[53],b[57],a[53]);
        
    
        and(andpr58[54],b[57],a[54]);
        
    
        and(andpr58[55],b[57],a[55]);
        
    
        and(andpr58[56],b[57],a[56]);
        
    
        and(andpr58[57],b[57],a[57]);
        
    
        and(andpr58[58],b[57],a[58]);
        
    
        and(andpr58[59],b[57],a[59]);
        
    
        and(andpr58[60],b[57],a[60]);
        
    
        and(andpr58[61],b[57],a[61]);
        
    
        and(andpr58[62],b[57],a[62]);
        
    
        and(andpr58[63],b[57],a[63]);
        
    
    not(si[57],andpr58[63]);

    
        and(andpr59[0],b[58],a[0]);
        
    
        and(andpr59[1],b[58],a[1]);
        
    
        and(andpr59[2],b[58],a[2]);
        
    
        and(andpr59[3],b[58],a[3]);
        
    
        and(andpr59[4],b[58],a[4]);
        
    
        and(andpr59[5],b[58],a[5]);
        
    
        and(andpr59[6],b[58],a[6]);
        
    
        and(andpr59[7],b[58],a[7]);
        
    
        and(andpr59[8],b[58],a[8]);
        
    
        and(andpr59[9],b[58],a[9]);
        
    
        and(andpr59[10],b[58],a[10]);
        
    
        and(andpr59[11],b[58],a[11]);
        
    
        and(andpr59[12],b[58],a[12]);
        
    
        and(andpr59[13],b[58],a[13]);
        
    
        and(andpr59[14],b[58],a[14]);
        
    
        and(andpr59[15],b[58],a[15]);
        
    
        and(andpr59[16],b[58],a[16]);
        
    
        and(andpr59[17],b[58],a[17]);
        
    
        and(andpr59[18],b[58],a[18]);
        
    
        and(andpr59[19],b[58],a[19]);
        
    
        and(andpr59[20],b[58],a[20]);
        
    
        and(andpr59[21],b[58],a[21]);
        
    
        and(andpr59[22],b[58],a[22]);
        
    
        and(andpr59[23],b[58],a[23]);
        
    
        and(andpr59[24],b[58],a[24]);
        
    
        and(andpr59[25],b[58],a[25]);
        
    
        and(andpr59[26],b[58],a[26]);
        
    
        and(andpr59[27],b[58],a[27]);
        
    
        and(andpr59[28],b[58],a[28]);
        
    
        and(andpr59[29],b[58],a[29]);
        
    
        and(andpr59[30],b[58],a[30]);
        
    
        and(andpr59[31],b[58],a[31]);
        
    
        and(andpr59[32],b[58],a[32]);
        
    
        and(andpr59[33],b[58],a[33]);
        
    
        and(andpr59[34],b[58],a[34]);
        
    
        and(andpr59[35],b[58],a[35]);
        
    
        and(andpr59[36],b[58],a[36]);
        
    
        and(andpr59[37],b[58],a[37]);
        
    
        and(andpr59[38],b[58],a[38]);
        
    
        and(andpr59[39],b[58],a[39]);
        
    
        and(andpr59[40],b[58],a[40]);
        
    
        and(andpr59[41],b[58],a[41]);
        
    
        and(andpr59[42],b[58],a[42]);
        
    
        and(andpr59[43],b[58],a[43]);
        
    
        and(andpr59[44],b[58],a[44]);
        
    
        and(andpr59[45],b[58],a[45]);
        
    
        and(andpr59[46],b[58],a[46]);
        
    
        and(andpr59[47],b[58],a[47]);
        
    
        and(andpr59[48],b[58],a[48]);
        
    
        and(andpr59[49],b[58],a[49]);
        
    
        and(andpr59[50],b[58],a[50]);
        
    
        and(andpr59[51],b[58],a[51]);
        
    
        and(andpr59[52],b[58],a[52]);
        
    
        and(andpr59[53],b[58],a[53]);
        
    
        and(andpr59[54],b[58],a[54]);
        
    
        and(andpr59[55],b[58],a[55]);
        
    
        and(andpr59[56],b[58],a[56]);
        
    
        and(andpr59[57],b[58],a[57]);
        
    
        and(andpr59[58],b[58],a[58]);
        
    
        and(andpr59[59],b[58],a[59]);
        
    
        and(andpr59[60],b[58],a[60]);
        
    
        and(andpr59[61],b[58],a[61]);
        
    
        and(andpr59[62],b[58],a[62]);
        
    
        and(andpr59[63],b[58],a[63]);
        
    
    not(si[58],andpr59[63]);

    
        and(andpr60[0],b[59],a[0]);
        
    
        and(andpr60[1],b[59],a[1]);
        
    
        and(andpr60[2],b[59],a[2]);
        
    
        and(andpr60[3],b[59],a[3]);
        
    
        and(andpr60[4],b[59],a[4]);
        
    
        and(andpr60[5],b[59],a[5]);
        
    
        and(andpr60[6],b[59],a[6]);
        
    
        and(andpr60[7],b[59],a[7]);
        
    
        and(andpr60[8],b[59],a[8]);
        
    
        and(andpr60[9],b[59],a[9]);
        
    
        and(andpr60[10],b[59],a[10]);
        
    
        and(andpr60[11],b[59],a[11]);
        
    
        and(andpr60[12],b[59],a[12]);
        
    
        and(andpr60[13],b[59],a[13]);
        
    
        and(andpr60[14],b[59],a[14]);
        
    
        and(andpr60[15],b[59],a[15]);
        
    
        and(andpr60[16],b[59],a[16]);
        
    
        and(andpr60[17],b[59],a[17]);
        
    
        and(andpr60[18],b[59],a[18]);
        
    
        and(andpr60[19],b[59],a[19]);
        
    
        and(andpr60[20],b[59],a[20]);
        
    
        and(andpr60[21],b[59],a[21]);
        
    
        and(andpr60[22],b[59],a[22]);
        
    
        and(andpr60[23],b[59],a[23]);
        
    
        and(andpr60[24],b[59],a[24]);
        
    
        and(andpr60[25],b[59],a[25]);
        
    
        and(andpr60[26],b[59],a[26]);
        
    
        and(andpr60[27],b[59],a[27]);
        
    
        and(andpr60[28],b[59],a[28]);
        
    
        and(andpr60[29],b[59],a[29]);
        
    
        and(andpr60[30],b[59],a[30]);
        
    
        and(andpr60[31],b[59],a[31]);
        
    
        and(andpr60[32],b[59],a[32]);
        
    
        and(andpr60[33],b[59],a[33]);
        
    
        and(andpr60[34],b[59],a[34]);
        
    
        and(andpr60[35],b[59],a[35]);
        
    
        and(andpr60[36],b[59],a[36]);
        
    
        and(andpr60[37],b[59],a[37]);
        
    
        and(andpr60[38],b[59],a[38]);
        
    
        and(andpr60[39],b[59],a[39]);
        
    
        and(andpr60[40],b[59],a[40]);
        
    
        and(andpr60[41],b[59],a[41]);
        
    
        and(andpr60[42],b[59],a[42]);
        
    
        and(andpr60[43],b[59],a[43]);
        
    
        and(andpr60[44],b[59],a[44]);
        
    
        and(andpr60[45],b[59],a[45]);
        
    
        and(andpr60[46],b[59],a[46]);
        
    
        and(andpr60[47],b[59],a[47]);
        
    
        and(andpr60[48],b[59],a[48]);
        
    
        and(andpr60[49],b[59],a[49]);
        
    
        and(andpr60[50],b[59],a[50]);
        
    
        and(andpr60[51],b[59],a[51]);
        
    
        and(andpr60[52],b[59],a[52]);
        
    
        and(andpr60[53],b[59],a[53]);
        
    
        and(andpr60[54],b[59],a[54]);
        
    
        and(andpr60[55],b[59],a[55]);
        
    
        and(andpr60[56],b[59],a[56]);
        
    
        and(andpr60[57],b[59],a[57]);
        
    
        and(andpr60[58],b[59],a[58]);
        
    
        and(andpr60[59],b[59],a[59]);
        
    
        and(andpr60[60],b[59],a[60]);
        
    
        and(andpr60[61],b[59],a[61]);
        
    
        and(andpr60[62],b[59],a[62]);
        
    
        and(andpr60[63],b[59],a[63]);
        
    
    not(si[59],andpr60[63]);

    
        and(andpr61[0],b[60],a[0]);
        
    
        and(andpr61[1],b[60],a[1]);
        
    
        and(andpr61[2],b[60],a[2]);
        
    
        and(andpr61[3],b[60],a[3]);
        
    
        and(andpr61[4],b[60],a[4]);
        
    
        and(andpr61[5],b[60],a[5]);
        
    
        and(andpr61[6],b[60],a[6]);
        
    
        and(andpr61[7],b[60],a[7]);
        
    
        and(andpr61[8],b[60],a[8]);
        
    
        and(andpr61[9],b[60],a[9]);
        
    
        and(andpr61[10],b[60],a[10]);
        
    
        and(andpr61[11],b[60],a[11]);
        
    
        and(andpr61[12],b[60],a[12]);
        
    
        and(andpr61[13],b[60],a[13]);
        
    
        and(andpr61[14],b[60],a[14]);
        
    
        and(andpr61[15],b[60],a[15]);
        
    
        and(andpr61[16],b[60],a[16]);
        
    
        and(andpr61[17],b[60],a[17]);
        
    
        and(andpr61[18],b[60],a[18]);
        
    
        and(andpr61[19],b[60],a[19]);
        
    
        and(andpr61[20],b[60],a[20]);
        
    
        and(andpr61[21],b[60],a[21]);
        
    
        and(andpr61[22],b[60],a[22]);
        
    
        and(andpr61[23],b[60],a[23]);
        
    
        and(andpr61[24],b[60],a[24]);
        
    
        and(andpr61[25],b[60],a[25]);
        
    
        and(andpr61[26],b[60],a[26]);
        
    
        and(andpr61[27],b[60],a[27]);
        
    
        and(andpr61[28],b[60],a[28]);
        
    
        and(andpr61[29],b[60],a[29]);
        
    
        and(andpr61[30],b[60],a[30]);
        
    
        and(andpr61[31],b[60],a[31]);
        
    
        and(andpr61[32],b[60],a[32]);
        
    
        and(andpr61[33],b[60],a[33]);
        
    
        and(andpr61[34],b[60],a[34]);
        
    
        and(andpr61[35],b[60],a[35]);
        
    
        and(andpr61[36],b[60],a[36]);
        
    
        and(andpr61[37],b[60],a[37]);
        
    
        and(andpr61[38],b[60],a[38]);
        
    
        and(andpr61[39],b[60],a[39]);
        
    
        and(andpr61[40],b[60],a[40]);
        
    
        and(andpr61[41],b[60],a[41]);
        
    
        and(andpr61[42],b[60],a[42]);
        
    
        and(andpr61[43],b[60],a[43]);
        
    
        and(andpr61[44],b[60],a[44]);
        
    
        and(andpr61[45],b[60],a[45]);
        
    
        and(andpr61[46],b[60],a[46]);
        
    
        and(andpr61[47],b[60],a[47]);
        
    
        and(andpr61[48],b[60],a[48]);
        
    
        and(andpr61[49],b[60],a[49]);
        
    
        and(andpr61[50],b[60],a[50]);
        
    
        and(andpr61[51],b[60],a[51]);
        
    
        and(andpr61[52],b[60],a[52]);
        
    
        and(andpr61[53],b[60],a[53]);
        
    
        and(andpr61[54],b[60],a[54]);
        
    
        and(andpr61[55],b[60],a[55]);
        
    
        and(andpr61[56],b[60],a[56]);
        
    
        and(andpr61[57],b[60],a[57]);
        
    
        and(andpr61[58],b[60],a[58]);
        
    
        and(andpr61[59],b[60],a[59]);
        
    
        and(andpr61[60],b[60],a[60]);
        
    
        and(andpr61[61],b[60],a[61]);
        
    
        and(andpr61[62],b[60],a[62]);
        
    
        and(andpr61[63],b[60],a[63]);
        
    
    not(si[60],andpr61[63]);

    
        and(andpr62[0],b[61],a[0]);
        
    
        and(andpr62[1],b[61],a[1]);
        
    
        and(andpr62[2],b[61],a[2]);
        
    
        and(andpr62[3],b[61],a[3]);
        
    
        and(andpr62[4],b[61],a[4]);
        
    
        and(andpr62[5],b[61],a[5]);
        
    
        and(andpr62[6],b[61],a[6]);
        
    
        and(andpr62[7],b[61],a[7]);
        
    
        and(andpr62[8],b[61],a[8]);
        
    
        and(andpr62[9],b[61],a[9]);
        
    
        and(andpr62[10],b[61],a[10]);
        
    
        and(andpr62[11],b[61],a[11]);
        
    
        and(andpr62[12],b[61],a[12]);
        
    
        and(andpr62[13],b[61],a[13]);
        
    
        and(andpr62[14],b[61],a[14]);
        
    
        and(andpr62[15],b[61],a[15]);
        
    
        and(andpr62[16],b[61],a[16]);
        
    
        and(andpr62[17],b[61],a[17]);
        
    
        and(andpr62[18],b[61],a[18]);
        
    
        and(andpr62[19],b[61],a[19]);
        
    
        and(andpr62[20],b[61],a[20]);
        
    
        and(andpr62[21],b[61],a[21]);
        
    
        and(andpr62[22],b[61],a[22]);
        
    
        and(andpr62[23],b[61],a[23]);
        
    
        and(andpr62[24],b[61],a[24]);
        
    
        and(andpr62[25],b[61],a[25]);
        
    
        and(andpr62[26],b[61],a[26]);
        
    
        and(andpr62[27],b[61],a[27]);
        
    
        and(andpr62[28],b[61],a[28]);
        
    
        and(andpr62[29],b[61],a[29]);
        
    
        and(andpr62[30],b[61],a[30]);
        
    
        and(andpr62[31],b[61],a[31]);
        
    
        and(andpr62[32],b[61],a[32]);
        
    
        and(andpr62[33],b[61],a[33]);
        
    
        and(andpr62[34],b[61],a[34]);
        
    
        and(andpr62[35],b[61],a[35]);
        
    
        and(andpr62[36],b[61],a[36]);
        
    
        and(andpr62[37],b[61],a[37]);
        
    
        and(andpr62[38],b[61],a[38]);
        
    
        and(andpr62[39],b[61],a[39]);
        
    
        and(andpr62[40],b[61],a[40]);
        
    
        and(andpr62[41],b[61],a[41]);
        
    
        and(andpr62[42],b[61],a[42]);
        
    
        and(andpr62[43],b[61],a[43]);
        
    
        and(andpr62[44],b[61],a[44]);
        
    
        and(andpr62[45],b[61],a[45]);
        
    
        and(andpr62[46],b[61],a[46]);
        
    
        and(andpr62[47],b[61],a[47]);
        
    
        and(andpr62[48],b[61],a[48]);
        
    
        and(andpr62[49],b[61],a[49]);
        
    
        and(andpr62[50],b[61],a[50]);
        
    
        and(andpr62[51],b[61],a[51]);
        
    
        and(andpr62[52],b[61],a[52]);
        
    
        and(andpr62[53],b[61],a[53]);
        
    
        and(andpr62[54],b[61],a[54]);
        
    
        and(andpr62[55],b[61],a[55]);
        
    
        and(andpr62[56],b[61],a[56]);
        
    
        and(andpr62[57],b[61],a[57]);
        
    
        and(andpr62[58],b[61],a[58]);
        
    
        and(andpr62[59],b[61],a[59]);
        
    
        and(andpr62[60],b[61],a[60]);
        
    
        and(andpr62[61],b[61],a[61]);
        
    
        and(andpr62[62],b[61],a[62]);
        
    
        and(andpr62[63],b[61],a[63]);
        
    
    not(si[61],andpr62[63]);

    
        and(andpr63[0],b[62],a[0]);
        
    
        and(andpr63[1],b[62],a[1]);
        
    
        and(andpr63[2],b[62],a[2]);
        
    
        and(andpr63[3],b[62],a[3]);
        
    
        and(andpr63[4],b[62],a[4]);
        
    
        and(andpr63[5],b[62],a[5]);
        
    
        and(andpr63[6],b[62],a[6]);
        
    
        and(andpr63[7],b[62],a[7]);
        
    
        and(andpr63[8],b[62],a[8]);
        
    
        and(andpr63[9],b[62],a[9]);
        
    
        and(andpr63[10],b[62],a[10]);
        
    
        and(andpr63[11],b[62],a[11]);
        
    
        and(andpr63[12],b[62],a[12]);
        
    
        and(andpr63[13],b[62],a[13]);
        
    
        and(andpr63[14],b[62],a[14]);
        
    
        and(andpr63[15],b[62],a[15]);
        
    
        and(andpr63[16],b[62],a[16]);
        
    
        and(andpr63[17],b[62],a[17]);
        
    
        and(andpr63[18],b[62],a[18]);
        
    
        and(andpr63[19],b[62],a[19]);
        
    
        and(andpr63[20],b[62],a[20]);
        
    
        and(andpr63[21],b[62],a[21]);
        
    
        and(andpr63[22],b[62],a[22]);
        
    
        and(andpr63[23],b[62],a[23]);
        
    
        and(andpr63[24],b[62],a[24]);
        
    
        and(andpr63[25],b[62],a[25]);
        
    
        and(andpr63[26],b[62],a[26]);
        
    
        and(andpr63[27],b[62],a[27]);
        
    
        and(andpr63[28],b[62],a[28]);
        
    
        and(andpr63[29],b[62],a[29]);
        
    
        and(andpr63[30],b[62],a[30]);
        
    
        and(andpr63[31],b[62],a[31]);
        
    
        and(andpr63[32],b[62],a[32]);
        
    
        and(andpr63[33],b[62],a[33]);
        
    
        and(andpr63[34],b[62],a[34]);
        
    
        and(andpr63[35],b[62],a[35]);
        
    
        and(andpr63[36],b[62],a[36]);
        
    
        and(andpr63[37],b[62],a[37]);
        
    
        and(andpr63[38],b[62],a[38]);
        
    
        and(andpr63[39],b[62],a[39]);
        
    
        and(andpr63[40],b[62],a[40]);
        
    
        and(andpr63[41],b[62],a[41]);
        
    
        and(andpr63[42],b[62],a[42]);
        
    
        and(andpr63[43],b[62],a[43]);
        
    
        and(andpr63[44],b[62],a[44]);
        
    
        and(andpr63[45],b[62],a[45]);
        
    
        and(andpr63[46],b[62],a[46]);
        
    
        and(andpr63[47],b[62],a[47]);
        
    
        and(andpr63[48],b[62],a[48]);
        
    
        and(andpr63[49],b[62],a[49]);
        
    
        and(andpr63[50],b[62],a[50]);
        
    
        and(andpr63[51],b[62],a[51]);
        
    
        and(andpr63[52],b[62],a[52]);
        
    
        and(andpr63[53],b[62],a[53]);
        
    
        and(andpr63[54],b[62],a[54]);
        
    
        and(andpr63[55],b[62],a[55]);
        
    
        and(andpr63[56],b[62],a[56]);
        
    
        and(andpr63[57],b[62],a[57]);
        
    
        and(andpr63[58],b[62],a[58]);
        
    
        and(andpr63[59],b[62],a[59]);
        
    
        and(andpr63[60],b[62],a[60]);
        
    
        and(andpr63[61],b[62],a[61]);
        
    
        and(andpr63[62],b[62],a[62]);
        
    
        and(andpr63[63],b[62],a[63]);
        
    
    not(si[62],andpr63[63]);


    and(andpr64[0],b[63],~a[0]);

    and(andpr64[1],b[63],~a[1]);

    and(andpr64[2],b[63],~a[2]);

    and(andpr64[3],b[63],~a[3]);

    and(andpr64[4],b[63],~a[4]);

    and(andpr64[5],b[63],~a[5]);

    and(andpr64[6],b[63],~a[6]);

    and(andpr64[7],b[63],~a[7]);

    and(andpr64[8],b[63],~a[8]);

    and(andpr64[9],b[63],~a[9]);

    and(andpr64[10],b[63],~a[10]);

    and(andpr64[11],b[63],~a[11]);

    and(andpr64[12],b[63],~a[12]);

    and(andpr64[13],b[63],~a[13]);

    and(andpr64[14],b[63],~a[14]);

    and(andpr64[15],b[63],~a[15]);

    and(andpr64[16],b[63],~a[16]);

    and(andpr64[17],b[63],~a[17]);

    and(andpr64[18],b[63],~a[18]);

    and(andpr64[19],b[63],~a[19]);

    and(andpr64[20],b[63],~a[20]);

    and(andpr64[21],b[63],~a[21]);

    and(andpr64[22],b[63],~a[22]);

    and(andpr64[23],b[63],~a[23]);

    and(andpr64[24],b[63],~a[24]);

    and(andpr64[25],b[63],~a[25]);

    and(andpr64[26],b[63],~a[26]);

    and(andpr64[27],b[63],~a[27]);

    and(andpr64[28],b[63],~a[28]);

    and(andpr64[29],b[63],~a[29]);

    and(andpr64[30],b[63],~a[30]);

    and(andpr64[31],b[63],~a[31]);

    and(andpr64[32],b[63],~a[32]);

    and(andpr64[33],b[63],~a[33]);

    and(andpr64[34],b[63],~a[34]);

    and(andpr64[35],b[63],~a[35]);

    and(andpr64[36],b[63],~a[36]);

    and(andpr64[37],b[63],~a[37]);

    and(andpr64[38],b[63],~a[38]);

    and(andpr64[39],b[63],~a[39]);

    and(andpr64[40],b[63],~a[40]);

    and(andpr64[41],b[63],~a[41]);

    and(andpr64[42],b[63],~a[42]);

    and(andpr64[43],b[63],~a[43]);

    and(andpr64[44],b[63],~a[44]);

    and(andpr64[45],b[63],~a[45]);

    and(andpr64[46],b[63],~a[46]);

    and(andpr64[47],b[63],~a[47]);

    and(andpr64[48],b[63],~a[48]);

    and(andpr64[49],b[63],~a[49]);

    and(andpr64[50],b[63],~a[50]);

    and(andpr64[51],b[63],~a[51]);

    and(andpr64[52],b[63],~a[52]);

    and(andpr64[53],b[63],~a[53]);

    and(andpr64[54],b[63],~a[54]);

    and(andpr64[55],b[63],~a[55]);

    and(andpr64[56],b[63],~a[56]);

    and(andpr64[57],b[63],~a[57]);

    and(andpr64[58],b[63],~a[58]);

    and(andpr64[59],b[63],~a[59]);

    and(andpr64[60],b[63],~a[60]);

    and(andpr64[61],b[63],~a[61]);

    and(andpr64[62],b[63],~a[62]);

    and(andpr64[63],b[63],~a[63]);

not(si[63],andpr64[63]);


half_adder ha1(andpr1[1],andpr2[0],c1[0],p[1]);


full_add fa1_1(andpr1[2],andpr2[1],andpr3[0],c1[1],s1[0]);


full_add fa1_2(andpr1[3],andpr2[2],andpr3[1],c1[2],s1[1]);


full_add fa1_3(andpr1[4],andpr2[3],andpr3[2],c1[3],s1[2]);


full_add fa1_4(andpr1[5],andpr2[4],andpr3[3],c1[4],s1[3]);


full_add fa1_5(andpr1[6],andpr2[5],andpr3[4],c1[5],s1[4]);


full_add fa1_6(andpr1[7],andpr2[6],andpr3[5],c1[6],s1[5]);


full_add fa1_7(andpr1[8],andpr2[7],andpr3[6],c1[7],s1[6]);


full_add fa1_8(andpr1[9],andpr2[8],andpr3[7],c1[8],s1[7]);


full_add fa1_9(andpr1[10],andpr2[9],andpr3[8],c1[9],s1[8]);


full_add fa1_10(andpr1[11],andpr2[10],andpr3[9],c1[10],s1[9]);


full_add fa1_11(andpr1[12],andpr2[11],andpr3[10],c1[11],s1[10]);


full_add fa1_12(andpr1[13],andpr2[12],andpr3[11],c1[12],s1[11]);


full_add fa1_13(andpr1[14],andpr2[13],andpr3[12],c1[13],s1[12]);


full_add fa1_14(andpr1[15],andpr2[14],andpr3[13],c1[14],s1[13]);


full_add fa1_15(andpr1[16],andpr2[15],andpr3[14],c1[15],s1[14]);


full_add fa1_16(andpr1[17],andpr2[16],andpr3[15],c1[16],s1[15]);


full_add fa1_17(andpr1[18],andpr2[17],andpr3[16],c1[17],s1[16]);


full_add fa1_18(andpr1[19],andpr2[18],andpr3[17],c1[18],s1[17]);


full_add fa1_19(andpr1[20],andpr2[19],andpr3[18],c1[19],s1[18]);


full_add fa1_20(andpr1[21],andpr2[20],andpr3[19],c1[20],s1[19]);


full_add fa1_21(andpr1[22],andpr2[21],andpr3[20],c1[21],s1[20]);


full_add fa1_22(andpr1[23],andpr2[22],andpr3[21],c1[22],s1[21]);


full_add fa1_23(andpr1[24],andpr2[23],andpr3[22],c1[23],s1[22]);


full_add fa1_24(andpr1[25],andpr2[24],andpr3[23],c1[24],s1[23]);


full_add fa1_25(andpr1[26],andpr2[25],andpr3[24],c1[25],s1[24]);


full_add fa1_26(andpr1[27],andpr2[26],andpr3[25],c1[26],s1[25]);


full_add fa1_27(andpr1[28],andpr2[27],andpr3[26],c1[27],s1[26]);


full_add fa1_28(andpr1[29],andpr2[28],andpr3[27],c1[28],s1[27]);


full_add fa1_29(andpr1[30],andpr2[29],andpr3[28],c1[29],s1[28]);


full_add fa1_30(andpr1[31],andpr2[30],andpr3[29],c1[30],s1[29]);


full_add fa1_31(andpr1[32],andpr2[31],andpr3[30],c1[31],s1[30]);


full_add fa1_32(andpr1[33],andpr2[32],andpr3[31],c1[32],s1[31]);


full_add fa1_33(andpr1[34],andpr2[33],andpr3[32],c1[33],s1[32]);


full_add fa1_34(andpr1[35],andpr2[34],andpr3[33],c1[34],s1[33]);


full_add fa1_35(andpr1[36],andpr2[35],andpr3[34],c1[35],s1[34]);


full_add fa1_36(andpr1[37],andpr2[36],andpr3[35],c1[36],s1[35]);


full_add fa1_37(andpr1[38],andpr2[37],andpr3[36],c1[37],s1[36]);


full_add fa1_38(andpr1[39],andpr2[38],andpr3[37],c1[38],s1[37]);


full_add fa1_39(andpr1[40],andpr2[39],andpr3[38],c1[39],s1[38]);


full_add fa1_40(andpr1[41],andpr2[40],andpr3[39],c1[40],s1[39]);


full_add fa1_41(andpr1[42],andpr2[41],andpr3[40],c1[41],s1[40]);


full_add fa1_42(andpr1[43],andpr2[42],andpr3[41],c1[42],s1[41]);


full_add fa1_43(andpr1[44],andpr2[43],andpr3[42],c1[43],s1[42]);


full_add fa1_44(andpr1[45],andpr2[44],andpr3[43],c1[44],s1[43]);


full_add fa1_45(andpr1[46],andpr2[45],andpr3[44],c1[45],s1[44]);


full_add fa1_46(andpr1[47],andpr2[46],andpr3[45],c1[46],s1[45]);


full_add fa1_47(andpr1[48],andpr2[47],andpr3[46],c1[47],s1[46]);


full_add fa1_48(andpr1[49],andpr2[48],andpr3[47],c1[48],s1[47]);


full_add fa1_49(andpr1[50],andpr2[49],andpr3[48],c1[49],s1[48]);


full_add fa1_50(andpr1[51],andpr2[50],andpr3[49],c1[50],s1[49]);


full_add fa1_51(andpr1[52],andpr2[51],andpr3[50],c1[51],s1[50]);


full_add fa1_52(andpr1[53],andpr2[52],andpr3[51],c1[52],s1[51]);


full_add fa1_53(andpr1[54],andpr2[53],andpr3[52],c1[53],s1[52]);


full_add fa1_54(andpr1[55],andpr2[54],andpr3[53],c1[54],s1[53]);


full_add fa1_55(andpr1[56],andpr2[55],andpr3[54],c1[55],s1[54]);


full_add fa1_56(andpr1[57],andpr2[56],andpr3[55],c1[56],s1[55]);


full_add fa1_57(andpr1[58],andpr2[57],andpr3[56],c1[57],s1[56]);


full_add fa1_58(andpr1[59],andpr2[58],andpr3[57],c1[58],s1[57]);


full_add fa1_59(andpr1[60],andpr2[59],andpr3[58],c1[59],s1[58]);


full_add fa1_60(andpr1[61],andpr2[60],andpr3[59],c1[60],s1[59]);


full_add fa1_61(andpr1[62],andpr2[61],andpr3[60],c1[61],s1[60]);


full_add fa1_62(andpr1[63],andpr2[62],andpr3[61],c1[62],s1[61]);



full_add fa2_63(si[0],si[1],andpr3[62],c1[63],s1[62]);



half_adder ha2(s1[0],c1[0],c2[0],p[2]);


full_add fa2_0(s1[1],c1[1],andpr4[0],c2[1],s2[0]);


full_add fa2_1(s1[2],c1[2],andpr4[1],c2[2],s2[1]);


full_add fa2_2(s1[3],c1[3],andpr4[2],c2[3],s2[2]);


full_add fa2_3(s1[4],c1[4],andpr4[3],c2[4],s2[3]);


full_add fa2_4(s1[5],c1[5],andpr4[4],c2[5],s2[4]);


full_add fa2_5(s1[6],c1[6],andpr4[5],c2[6],s2[5]);


full_add fa2_6(s1[7],c1[7],andpr4[6],c2[7],s2[6]);


full_add fa2_7(s1[8],c1[8],andpr4[7],c2[8],s2[7]);


full_add fa2_8(s1[9],c1[9],andpr4[8],c2[9],s2[8]);


full_add fa2_9(s1[10],c1[10],andpr4[9],c2[10],s2[9]);


full_add fa2_10(s1[11],c1[11],andpr4[10],c2[11],s2[10]);


full_add fa2_11(s1[12],c1[12],andpr4[11],c2[12],s2[11]);


full_add fa2_12(s1[13],c1[13],andpr4[12],c2[13],s2[12]);


full_add fa2_13(s1[14],c1[14],andpr4[13],c2[14],s2[13]);


full_add fa2_14(s1[15],c1[15],andpr4[14],c2[15],s2[14]);


full_add fa2_15(s1[16],c1[16],andpr4[15],c2[16],s2[15]);


full_add fa2_16(s1[17],c1[17],andpr4[16],c2[17],s2[16]);


full_add fa2_17(s1[18],c1[18],andpr4[17],c2[18],s2[17]);


full_add fa2_18(s1[19],c1[19],andpr4[18],c2[19],s2[18]);


full_add fa2_19(s1[20],c1[20],andpr4[19],c2[20],s2[19]);


full_add fa2_20(s1[21],c1[21],andpr4[20],c2[21],s2[20]);


full_add fa2_21(s1[22],c1[22],andpr4[21],c2[22],s2[21]);


full_add fa2_22(s1[23],c1[23],andpr4[22],c2[23],s2[22]);


full_add fa2_23(s1[24],c1[24],andpr4[23],c2[24],s2[23]);


full_add fa2_24(s1[25],c1[25],andpr4[24],c2[25],s2[24]);


full_add fa2_25(s1[26],c1[26],andpr4[25],c2[26],s2[25]);


full_add fa2_26(s1[27],c1[27],andpr4[26],c2[27],s2[26]);


full_add fa2_27(s1[28],c1[28],andpr4[27],c2[28],s2[27]);


full_add fa2_28(s1[29],c1[29],andpr4[28],c2[29],s2[28]);


full_add fa2_29(s1[30],c1[30],andpr4[29],c2[30],s2[29]);


full_add fa2_30(s1[31],c1[31],andpr4[30],c2[31],s2[30]);


full_add fa2_31(s1[32],c1[32],andpr4[31],c2[32],s2[31]);


full_add fa2_32(s1[33],c1[33],andpr4[32],c2[33],s2[32]);


full_add fa2_33(s1[34],c1[34],andpr4[33],c2[34],s2[33]);


full_add fa2_34(s1[35],c1[35],andpr4[34],c2[35],s2[34]);


full_add fa2_35(s1[36],c1[36],andpr4[35],c2[36],s2[35]);


full_add fa2_36(s1[37],c1[37],andpr4[36],c2[37],s2[36]);


full_add fa2_37(s1[38],c1[38],andpr4[37],c2[38],s2[37]);


full_add fa2_38(s1[39],c1[39],andpr4[38],c2[39],s2[38]);


full_add fa2_39(s1[40],c1[40],andpr4[39],c2[40],s2[39]);


full_add fa2_40(s1[41],c1[41],andpr4[40],c2[41],s2[40]);


full_add fa2_41(s1[42],c1[42],andpr4[41],c2[42],s2[41]);


full_add fa2_42(s1[43],c1[43],andpr4[42],c2[43],s2[42]);


full_add fa2_43(s1[44],c1[44],andpr4[43],c2[44],s2[43]);


full_add fa2_44(s1[45],c1[45],andpr4[44],c2[45],s2[44]);


full_add fa2_45(s1[46],c1[46],andpr4[45],c2[46],s2[45]);


full_add fa2_46(s1[47],c1[47],andpr4[46],c2[47],s2[46]);


full_add fa2_47(s1[48],c1[48],andpr4[47],c2[48],s2[47]);


full_add fa2_48(s1[49],c1[49],andpr4[48],c2[49],s2[48]);


full_add fa2_49(s1[50],c1[50],andpr4[49],c2[50],s2[49]);


full_add fa2_50(s1[51],c1[51],andpr4[50],c2[51],s2[50]);


full_add fa2_51(s1[52],c1[52],andpr4[51],c2[52],s2[51]);


full_add fa2_52(s1[53],c1[53],andpr4[52],c2[53],s2[52]);


full_add fa2_53(s1[54],c1[54],andpr4[53],c2[54],s2[53]);


full_add fa2_54(s1[55],c1[55],andpr4[54],c2[55],s2[54]);


full_add fa2_55(s1[56],c1[56],andpr4[55],c2[56],s2[55]);


full_add fa2_56(s1[57],c1[57],andpr4[56],c2[57],s2[56]);


full_add fa2_57(s1[58],c1[58],andpr4[57],c2[58],s2[57]);


full_add fa2_58(s1[59],c1[59],andpr4[58],c2[59],s2[58]);


full_add fa2_59(s1[60],c1[60],andpr4[59],c2[60],s2[59]);


full_add fa2_60(s1[61],c1[61],andpr4[60],c2[61],s2[60]);


full_add fa2_61(s1[62],c1[62],andpr4[61],c2[62],s2[61]);


full_add fa2_62(si[2],c1[63],andpr4[62],c2[63],s2[62]);



half_adder ha3(s2[0],c2[0],c3[0],p[3]);


full_add fa3_0(s2[1],c2[1],andpr5[0],c3[1],s3[0]);


full_add fa3_1(s2[2],c2[2],andpr5[1],c3[2],s3[1]);


full_add fa3_2(s2[3],c2[3],andpr5[2],c3[3],s3[2]);


full_add fa3_3(s2[4],c2[4],andpr5[3],c3[4],s3[3]);


full_add fa3_4(s2[5],c2[5],andpr5[4],c3[5],s3[4]);


full_add fa3_5(s2[6],c2[6],andpr5[5],c3[6],s3[5]);


full_add fa3_6(s2[7],c2[7],andpr5[6],c3[7],s3[6]);


full_add fa3_7(s2[8],c2[8],andpr5[7],c3[8],s3[7]);


full_add fa3_8(s2[9],c2[9],andpr5[8],c3[9],s3[8]);


full_add fa3_9(s2[10],c2[10],andpr5[9],c3[10],s3[9]);


full_add fa3_10(s2[11],c2[11],andpr5[10],c3[11],s3[10]);


full_add fa3_11(s2[12],c2[12],andpr5[11],c3[12],s3[11]);


full_add fa3_12(s2[13],c2[13],andpr5[12],c3[13],s3[12]);


full_add fa3_13(s2[14],c2[14],andpr5[13],c3[14],s3[13]);


full_add fa3_14(s2[15],c2[15],andpr5[14],c3[15],s3[14]);


full_add fa3_15(s2[16],c2[16],andpr5[15],c3[16],s3[15]);


full_add fa3_16(s2[17],c2[17],andpr5[16],c3[17],s3[16]);


full_add fa3_17(s2[18],c2[18],andpr5[17],c3[18],s3[17]);


full_add fa3_18(s2[19],c2[19],andpr5[18],c3[19],s3[18]);


full_add fa3_19(s2[20],c2[20],andpr5[19],c3[20],s3[19]);


full_add fa3_20(s2[21],c2[21],andpr5[20],c3[21],s3[20]);


full_add fa3_21(s2[22],c2[22],andpr5[21],c3[22],s3[21]);


full_add fa3_22(s2[23],c2[23],andpr5[22],c3[23],s3[22]);


full_add fa3_23(s2[24],c2[24],andpr5[23],c3[24],s3[23]);


full_add fa3_24(s2[25],c2[25],andpr5[24],c3[25],s3[24]);


full_add fa3_25(s2[26],c2[26],andpr5[25],c3[26],s3[25]);


full_add fa3_26(s2[27],c2[27],andpr5[26],c3[27],s3[26]);


full_add fa3_27(s2[28],c2[28],andpr5[27],c3[28],s3[27]);


full_add fa3_28(s2[29],c2[29],andpr5[28],c3[29],s3[28]);


full_add fa3_29(s2[30],c2[30],andpr5[29],c3[30],s3[29]);


full_add fa3_30(s2[31],c2[31],andpr5[30],c3[31],s3[30]);


full_add fa3_31(s2[32],c2[32],andpr5[31],c3[32],s3[31]);


full_add fa3_32(s2[33],c2[33],andpr5[32],c3[33],s3[32]);


full_add fa3_33(s2[34],c2[34],andpr5[33],c3[34],s3[33]);


full_add fa3_34(s2[35],c2[35],andpr5[34],c3[35],s3[34]);


full_add fa3_35(s2[36],c2[36],andpr5[35],c3[36],s3[35]);


full_add fa3_36(s2[37],c2[37],andpr5[36],c3[37],s3[36]);


full_add fa3_37(s2[38],c2[38],andpr5[37],c3[38],s3[37]);


full_add fa3_38(s2[39],c2[39],andpr5[38],c3[39],s3[38]);


full_add fa3_39(s2[40],c2[40],andpr5[39],c3[40],s3[39]);


full_add fa3_40(s2[41],c2[41],andpr5[40],c3[41],s3[40]);


full_add fa3_41(s2[42],c2[42],andpr5[41],c3[42],s3[41]);


full_add fa3_42(s2[43],c2[43],andpr5[42],c3[43],s3[42]);


full_add fa3_43(s2[44],c2[44],andpr5[43],c3[44],s3[43]);


full_add fa3_44(s2[45],c2[45],andpr5[44],c3[45],s3[44]);


full_add fa3_45(s2[46],c2[46],andpr5[45],c3[46],s3[45]);


full_add fa3_46(s2[47],c2[47],andpr5[46],c3[47],s3[46]);


full_add fa3_47(s2[48],c2[48],andpr5[47],c3[48],s3[47]);


full_add fa3_48(s2[49],c2[49],andpr5[48],c3[49],s3[48]);


full_add fa3_49(s2[50],c2[50],andpr5[49],c3[50],s3[49]);


full_add fa3_50(s2[51],c2[51],andpr5[50],c3[51],s3[50]);


full_add fa3_51(s2[52],c2[52],andpr5[51],c3[52],s3[51]);


full_add fa3_52(s2[53],c2[53],andpr5[52],c3[53],s3[52]);


full_add fa3_53(s2[54],c2[54],andpr5[53],c3[54],s3[53]);


full_add fa3_54(s2[55],c2[55],andpr5[54],c3[55],s3[54]);


full_add fa3_55(s2[56],c2[56],andpr5[55],c3[56],s3[55]);


full_add fa3_56(s2[57],c2[57],andpr5[56],c3[57],s3[56]);


full_add fa3_57(s2[58],c2[58],andpr5[57],c3[58],s3[57]);


full_add fa3_58(s2[59],c2[59],andpr5[58],c3[59],s3[58]);


full_add fa3_59(s2[60],c2[60],andpr5[59],c3[60],s3[59]);


full_add fa3_60(s2[61],c2[61],andpr5[60],c3[61],s3[60]);


full_add fa3_61(s2[62],c2[62],andpr5[61],c3[62],s3[61]);


full_add fa3_62(si[3],c2[63],andpr5[62],c3[63],s3[62]);



half_adder ha4(s3[0],c3[0],c4[0],p[4]);


full_add fa4_0(s3[1],c3[1],andpr6[0],c4[1],s4[0]);


full_add fa4_1(s3[2],c3[2],andpr6[1],c4[2],s4[1]);


full_add fa4_2(s3[3],c3[3],andpr6[2],c4[3],s4[2]);


full_add fa4_3(s3[4],c3[4],andpr6[3],c4[4],s4[3]);


full_add fa4_4(s3[5],c3[5],andpr6[4],c4[5],s4[4]);


full_add fa4_5(s3[6],c3[6],andpr6[5],c4[6],s4[5]);


full_add fa4_6(s3[7],c3[7],andpr6[6],c4[7],s4[6]);


full_add fa4_7(s3[8],c3[8],andpr6[7],c4[8],s4[7]);


full_add fa4_8(s3[9],c3[9],andpr6[8],c4[9],s4[8]);


full_add fa4_9(s3[10],c3[10],andpr6[9],c4[10],s4[9]);


full_add fa4_10(s3[11],c3[11],andpr6[10],c4[11],s4[10]);


full_add fa4_11(s3[12],c3[12],andpr6[11],c4[12],s4[11]);


full_add fa4_12(s3[13],c3[13],andpr6[12],c4[13],s4[12]);


full_add fa4_13(s3[14],c3[14],andpr6[13],c4[14],s4[13]);


full_add fa4_14(s3[15],c3[15],andpr6[14],c4[15],s4[14]);


full_add fa4_15(s3[16],c3[16],andpr6[15],c4[16],s4[15]);


full_add fa4_16(s3[17],c3[17],andpr6[16],c4[17],s4[16]);


full_add fa4_17(s3[18],c3[18],andpr6[17],c4[18],s4[17]);


full_add fa4_18(s3[19],c3[19],andpr6[18],c4[19],s4[18]);


full_add fa4_19(s3[20],c3[20],andpr6[19],c4[20],s4[19]);


full_add fa4_20(s3[21],c3[21],andpr6[20],c4[21],s4[20]);


full_add fa4_21(s3[22],c3[22],andpr6[21],c4[22],s4[21]);


full_add fa4_22(s3[23],c3[23],andpr6[22],c4[23],s4[22]);


full_add fa4_23(s3[24],c3[24],andpr6[23],c4[24],s4[23]);


full_add fa4_24(s3[25],c3[25],andpr6[24],c4[25],s4[24]);


full_add fa4_25(s3[26],c3[26],andpr6[25],c4[26],s4[25]);


full_add fa4_26(s3[27],c3[27],andpr6[26],c4[27],s4[26]);


full_add fa4_27(s3[28],c3[28],andpr6[27],c4[28],s4[27]);


full_add fa4_28(s3[29],c3[29],andpr6[28],c4[29],s4[28]);


full_add fa4_29(s3[30],c3[30],andpr6[29],c4[30],s4[29]);


full_add fa4_30(s3[31],c3[31],andpr6[30],c4[31],s4[30]);


full_add fa4_31(s3[32],c3[32],andpr6[31],c4[32],s4[31]);


full_add fa4_32(s3[33],c3[33],andpr6[32],c4[33],s4[32]);


full_add fa4_33(s3[34],c3[34],andpr6[33],c4[34],s4[33]);


full_add fa4_34(s3[35],c3[35],andpr6[34],c4[35],s4[34]);


full_add fa4_35(s3[36],c3[36],andpr6[35],c4[36],s4[35]);


full_add fa4_36(s3[37],c3[37],andpr6[36],c4[37],s4[36]);


full_add fa4_37(s3[38],c3[38],andpr6[37],c4[38],s4[37]);


full_add fa4_38(s3[39],c3[39],andpr6[38],c4[39],s4[38]);


full_add fa4_39(s3[40],c3[40],andpr6[39],c4[40],s4[39]);


full_add fa4_40(s3[41],c3[41],andpr6[40],c4[41],s4[40]);


full_add fa4_41(s3[42],c3[42],andpr6[41],c4[42],s4[41]);


full_add fa4_42(s3[43],c3[43],andpr6[42],c4[43],s4[42]);


full_add fa4_43(s3[44],c3[44],andpr6[43],c4[44],s4[43]);


full_add fa4_44(s3[45],c3[45],andpr6[44],c4[45],s4[44]);


full_add fa4_45(s3[46],c3[46],andpr6[45],c4[46],s4[45]);


full_add fa4_46(s3[47],c3[47],andpr6[46],c4[47],s4[46]);


full_add fa4_47(s3[48],c3[48],andpr6[47],c4[48],s4[47]);


full_add fa4_48(s3[49],c3[49],andpr6[48],c4[49],s4[48]);


full_add fa4_49(s3[50],c3[50],andpr6[49],c4[50],s4[49]);


full_add fa4_50(s3[51],c3[51],andpr6[50],c4[51],s4[50]);


full_add fa4_51(s3[52],c3[52],andpr6[51],c4[52],s4[51]);


full_add fa4_52(s3[53],c3[53],andpr6[52],c4[53],s4[52]);


full_add fa4_53(s3[54],c3[54],andpr6[53],c4[54],s4[53]);


full_add fa4_54(s3[55],c3[55],andpr6[54],c4[55],s4[54]);


full_add fa4_55(s3[56],c3[56],andpr6[55],c4[56],s4[55]);


full_add fa4_56(s3[57],c3[57],andpr6[56],c4[57],s4[56]);


full_add fa4_57(s3[58],c3[58],andpr6[57],c4[58],s4[57]);


full_add fa4_58(s3[59],c3[59],andpr6[58],c4[59],s4[58]);


full_add fa4_59(s3[60],c3[60],andpr6[59],c4[60],s4[59]);


full_add fa4_60(s3[61],c3[61],andpr6[60],c4[61],s4[60]);


full_add fa4_61(s3[62],c3[62],andpr6[61],c4[62],s4[61]);


full_add fa4_62(si[4],c3[63],andpr6[62],c4[63],s4[62]);



half_adder ha5(s4[0],c4[0],c5[0],p[5]);


full_add fa5_0(s4[1],c4[1],andpr7[0],c5[1],s5[0]);


full_add fa5_1(s4[2],c4[2],andpr7[1],c5[2],s5[1]);


full_add fa5_2(s4[3],c4[3],andpr7[2],c5[3],s5[2]);


full_add fa5_3(s4[4],c4[4],andpr7[3],c5[4],s5[3]);


full_add fa5_4(s4[5],c4[5],andpr7[4],c5[5],s5[4]);


full_add fa5_5(s4[6],c4[6],andpr7[5],c5[6],s5[5]);


full_add fa5_6(s4[7],c4[7],andpr7[6],c5[7],s5[6]);


full_add fa5_7(s4[8],c4[8],andpr7[7],c5[8],s5[7]);


full_add fa5_8(s4[9],c4[9],andpr7[8],c5[9],s5[8]);


full_add fa5_9(s4[10],c4[10],andpr7[9],c5[10],s5[9]);


full_add fa5_10(s4[11],c4[11],andpr7[10],c5[11],s5[10]);


full_add fa5_11(s4[12],c4[12],andpr7[11],c5[12],s5[11]);


full_add fa5_12(s4[13],c4[13],andpr7[12],c5[13],s5[12]);


full_add fa5_13(s4[14],c4[14],andpr7[13],c5[14],s5[13]);


full_add fa5_14(s4[15],c4[15],andpr7[14],c5[15],s5[14]);


full_add fa5_15(s4[16],c4[16],andpr7[15],c5[16],s5[15]);


full_add fa5_16(s4[17],c4[17],andpr7[16],c5[17],s5[16]);


full_add fa5_17(s4[18],c4[18],andpr7[17],c5[18],s5[17]);


full_add fa5_18(s4[19],c4[19],andpr7[18],c5[19],s5[18]);


full_add fa5_19(s4[20],c4[20],andpr7[19],c5[20],s5[19]);


full_add fa5_20(s4[21],c4[21],andpr7[20],c5[21],s5[20]);


full_add fa5_21(s4[22],c4[22],andpr7[21],c5[22],s5[21]);


full_add fa5_22(s4[23],c4[23],andpr7[22],c5[23],s5[22]);


full_add fa5_23(s4[24],c4[24],andpr7[23],c5[24],s5[23]);


full_add fa5_24(s4[25],c4[25],andpr7[24],c5[25],s5[24]);


full_add fa5_25(s4[26],c4[26],andpr7[25],c5[26],s5[25]);


full_add fa5_26(s4[27],c4[27],andpr7[26],c5[27],s5[26]);


full_add fa5_27(s4[28],c4[28],andpr7[27],c5[28],s5[27]);


full_add fa5_28(s4[29],c4[29],andpr7[28],c5[29],s5[28]);


full_add fa5_29(s4[30],c4[30],andpr7[29],c5[30],s5[29]);


full_add fa5_30(s4[31],c4[31],andpr7[30],c5[31],s5[30]);


full_add fa5_31(s4[32],c4[32],andpr7[31],c5[32],s5[31]);


full_add fa5_32(s4[33],c4[33],andpr7[32],c5[33],s5[32]);


full_add fa5_33(s4[34],c4[34],andpr7[33],c5[34],s5[33]);


full_add fa5_34(s4[35],c4[35],andpr7[34],c5[35],s5[34]);


full_add fa5_35(s4[36],c4[36],andpr7[35],c5[36],s5[35]);


full_add fa5_36(s4[37],c4[37],andpr7[36],c5[37],s5[36]);


full_add fa5_37(s4[38],c4[38],andpr7[37],c5[38],s5[37]);


full_add fa5_38(s4[39],c4[39],andpr7[38],c5[39],s5[38]);


full_add fa5_39(s4[40],c4[40],andpr7[39],c5[40],s5[39]);


full_add fa5_40(s4[41],c4[41],andpr7[40],c5[41],s5[40]);


full_add fa5_41(s4[42],c4[42],andpr7[41],c5[42],s5[41]);


full_add fa5_42(s4[43],c4[43],andpr7[42],c5[43],s5[42]);


full_add fa5_43(s4[44],c4[44],andpr7[43],c5[44],s5[43]);


full_add fa5_44(s4[45],c4[45],andpr7[44],c5[45],s5[44]);


full_add fa5_45(s4[46],c4[46],andpr7[45],c5[46],s5[45]);


full_add fa5_46(s4[47],c4[47],andpr7[46],c5[47],s5[46]);


full_add fa5_47(s4[48],c4[48],andpr7[47],c5[48],s5[47]);


full_add fa5_48(s4[49],c4[49],andpr7[48],c5[49],s5[48]);


full_add fa5_49(s4[50],c4[50],andpr7[49],c5[50],s5[49]);


full_add fa5_50(s4[51],c4[51],andpr7[50],c5[51],s5[50]);


full_add fa5_51(s4[52],c4[52],andpr7[51],c5[52],s5[51]);


full_add fa5_52(s4[53],c4[53],andpr7[52],c5[53],s5[52]);


full_add fa5_53(s4[54],c4[54],andpr7[53],c5[54],s5[53]);


full_add fa5_54(s4[55],c4[55],andpr7[54],c5[55],s5[54]);


full_add fa5_55(s4[56],c4[56],andpr7[55],c5[56],s5[55]);


full_add fa5_56(s4[57],c4[57],andpr7[56],c5[57],s5[56]);


full_add fa5_57(s4[58],c4[58],andpr7[57],c5[58],s5[57]);


full_add fa5_58(s4[59],c4[59],andpr7[58],c5[59],s5[58]);


full_add fa5_59(s4[60],c4[60],andpr7[59],c5[60],s5[59]);


full_add fa5_60(s4[61],c4[61],andpr7[60],c5[61],s5[60]);


full_add fa5_61(s4[62],c4[62],andpr7[61],c5[62],s5[61]);


full_add fa5_62(si[5],c4[63],andpr7[62],c5[63],s5[62]);



half_adder ha6(s5[0],c5[0],c6[0],p[6]);


full_add fa6_0(s5[1],c5[1],andpr8[0],c6[1],s6[0]);


full_add fa6_1(s5[2],c5[2],andpr8[1],c6[2],s6[1]);


full_add fa6_2(s5[3],c5[3],andpr8[2],c6[3],s6[2]);


full_add fa6_3(s5[4],c5[4],andpr8[3],c6[4],s6[3]);


full_add fa6_4(s5[5],c5[5],andpr8[4],c6[5],s6[4]);


full_add fa6_5(s5[6],c5[6],andpr8[5],c6[6],s6[5]);


full_add fa6_6(s5[7],c5[7],andpr8[6],c6[7],s6[6]);


full_add fa6_7(s5[8],c5[8],andpr8[7],c6[8],s6[7]);


full_add fa6_8(s5[9],c5[9],andpr8[8],c6[9],s6[8]);


full_add fa6_9(s5[10],c5[10],andpr8[9],c6[10],s6[9]);


full_add fa6_10(s5[11],c5[11],andpr8[10],c6[11],s6[10]);


full_add fa6_11(s5[12],c5[12],andpr8[11],c6[12],s6[11]);


full_add fa6_12(s5[13],c5[13],andpr8[12],c6[13],s6[12]);


full_add fa6_13(s5[14],c5[14],andpr8[13],c6[14],s6[13]);


full_add fa6_14(s5[15],c5[15],andpr8[14],c6[15],s6[14]);


full_add fa6_15(s5[16],c5[16],andpr8[15],c6[16],s6[15]);


full_add fa6_16(s5[17],c5[17],andpr8[16],c6[17],s6[16]);


full_add fa6_17(s5[18],c5[18],andpr8[17],c6[18],s6[17]);


full_add fa6_18(s5[19],c5[19],andpr8[18],c6[19],s6[18]);


full_add fa6_19(s5[20],c5[20],andpr8[19],c6[20],s6[19]);


full_add fa6_20(s5[21],c5[21],andpr8[20],c6[21],s6[20]);


full_add fa6_21(s5[22],c5[22],andpr8[21],c6[22],s6[21]);


full_add fa6_22(s5[23],c5[23],andpr8[22],c6[23],s6[22]);


full_add fa6_23(s5[24],c5[24],andpr8[23],c6[24],s6[23]);


full_add fa6_24(s5[25],c5[25],andpr8[24],c6[25],s6[24]);


full_add fa6_25(s5[26],c5[26],andpr8[25],c6[26],s6[25]);


full_add fa6_26(s5[27],c5[27],andpr8[26],c6[27],s6[26]);


full_add fa6_27(s5[28],c5[28],andpr8[27],c6[28],s6[27]);


full_add fa6_28(s5[29],c5[29],andpr8[28],c6[29],s6[28]);


full_add fa6_29(s5[30],c5[30],andpr8[29],c6[30],s6[29]);


full_add fa6_30(s5[31],c5[31],andpr8[30],c6[31],s6[30]);


full_add fa6_31(s5[32],c5[32],andpr8[31],c6[32],s6[31]);


full_add fa6_32(s5[33],c5[33],andpr8[32],c6[33],s6[32]);


full_add fa6_33(s5[34],c5[34],andpr8[33],c6[34],s6[33]);


full_add fa6_34(s5[35],c5[35],andpr8[34],c6[35],s6[34]);


full_add fa6_35(s5[36],c5[36],andpr8[35],c6[36],s6[35]);


full_add fa6_36(s5[37],c5[37],andpr8[36],c6[37],s6[36]);


full_add fa6_37(s5[38],c5[38],andpr8[37],c6[38],s6[37]);


full_add fa6_38(s5[39],c5[39],andpr8[38],c6[39],s6[38]);


full_add fa6_39(s5[40],c5[40],andpr8[39],c6[40],s6[39]);


full_add fa6_40(s5[41],c5[41],andpr8[40],c6[41],s6[40]);


full_add fa6_41(s5[42],c5[42],andpr8[41],c6[42],s6[41]);


full_add fa6_42(s5[43],c5[43],andpr8[42],c6[43],s6[42]);


full_add fa6_43(s5[44],c5[44],andpr8[43],c6[44],s6[43]);


full_add fa6_44(s5[45],c5[45],andpr8[44],c6[45],s6[44]);


full_add fa6_45(s5[46],c5[46],andpr8[45],c6[46],s6[45]);


full_add fa6_46(s5[47],c5[47],andpr8[46],c6[47],s6[46]);


full_add fa6_47(s5[48],c5[48],andpr8[47],c6[48],s6[47]);


full_add fa6_48(s5[49],c5[49],andpr8[48],c6[49],s6[48]);


full_add fa6_49(s5[50],c5[50],andpr8[49],c6[50],s6[49]);


full_add fa6_50(s5[51],c5[51],andpr8[50],c6[51],s6[50]);


full_add fa6_51(s5[52],c5[52],andpr8[51],c6[52],s6[51]);


full_add fa6_52(s5[53],c5[53],andpr8[52],c6[53],s6[52]);


full_add fa6_53(s5[54],c5[54],andpr8[53],c6[54],s6[53]);


full_add fa6_54(s5[55],c5[55],andpr8[54],c6[55],s6[54]);


full_add fa6_55(s5[56],c5[56],andpr8[55],c6[56],s6[55]);


full_add fa6_56(s5[57],c5[57],andpr8[56],c6[57],s6[56]);


full_add fa6_57(s5[58],c5[58],andpr8[57],c6[58],s6[57]);


full_add fa6_58(s5[59],c5[59],andpr8[58],c6[59],s6[58]);


full_add fa6_59(s5[60],c5[60],andpr8[59],c6[60],s6[59]);


full_add fa6_60(s5[61],c5[61],andpr8[60],c6[61],s6[60]);


full_add fa6_61(s5[62],c5[62],andpr8[61],c6[62],s6[61]);


full_add fa6_62(si[6],c5[63],andpr8[62],c6[63],s6[62]);



half_adder ha7(s6[0],c6[0],c7[0],p[7]);


full_add fa7_0(s6[1],c6[1],andpr9[0],c7[1],s7[0]);


full_add fa7_1(s6[2],c6[2],andpr9[1],c7[2],s7[1]);


full_add fa7_2(s6[3],c6[3],andpr9[2],c7[3],s7[2]);


full_add fa7_3(s6[4],c6[4],andpr9[3],c7[4],s7[3]);


full_add fa7_4(s6[5],c6[5],andpr9[4],c7[5],s7[4]);


full_add fa7_5(s6[6],c6[6],andpr9[5],c7[6],s7[5]);


full_add fa7_6(s6[7],c6[7],andpr9[6],c7[7],s7[6]);


full_add fa7_7(s6[8],c6[8],andpr9[7],c7[8],s7[7]);


full_add fa7_8(s6[9],c6[9],andpr9[8],c7[9],s7[8]);


full_add fa7_9(s6[10],c6[10],andpr9[9],c7[10],s7[9]);


full_add fa7_10(s6[11],c6[11],andpr9[10],c7[11],s7[10]);


full_add fa7_11(s6[12],c6[12],andpr9[11],c7[12],s7[11]);


full_add fa7_12(s6[13],c6[13],andpr9[12],c7[13],s7[12]);


full_add fa7_13(s6[14],c6[14],andpr9[13],c7[14],s7[13]);


full_add fa7_14(s6[15],c6[15],andpr9[14],c7[15],s7[14]);


full_add fa7_15(s6[16],c6[16],andpr9[15],c7[16],s7[15]);


full_add fa7_16(s6[17],c6[17],andpr9[16],c7[17],s7[16]);


full_add fa7_17(s6[18],c6[18],andpr9[17],c7[18],s7[17]);


full_add fa7_18(s6[19],c6[19],andpr9[18],c7[19],s7[18]);


full_add fa7_19(s6[20],c6[20],andpr9[19],c7[20],s7[19]);


full_add fa7_20(s6[21],c6[21],andpr9[20],c7[21],s7[20]);


full_add fa7_21(s6[22],c6[22],andpr9[21],c7[22],s7[21]);


full_add fa7_22(s6[23],c6[23],andpr9[22],c7[23],s7[22]);


full_add fa7_23(s6[24],c6[24],andpr9[23],c7[24],s7[23]);


full_add fa7_24(s6[25],c6[25],andpr9[24],c7[25],s7[24]);


full_add fa7_25(s6[26],c6[26],andpr9[25],c7[26],s7[25]);


full_add fa7_26(s6[27],c6[27],andpr9[26],c7[27],s7[26]);


full_add fa7_27(s6[28],c6[28],andpr9[27],c7[28],s7[27]);


full_add fa7_28(s6[29],c6[29],andpr9[28],c7[29],s7[28]);


full_add fa7_29(s6[30],c6[30],andpr9[29],c7[30],s7[29]);


full_add fa7_30(s6[31],c6[31],andpr9[30],c7[31],s7[30]);


full_add fa7_31(s6[32],c6[32],andpr9[31],c7[32],s7[31]);


full_add fa7_32(s6[33],c6[33],andpr9[32],c7[33],s7[32]);


full_add fa7_33(s6[34],c6[34],andpr9[33],c7[34],s7[33]);


full_add fa7_34(s6[35],c6[35],andpr9[34],c7[35],s7[34]);


full_add fa7_35(s6[36],c6[36],andpr9[35],c7[36],s7[35]);


full_add fa7_36(s6[37],c6[37],andpr9[36],c7[37],s7[36]);


full_add fa7_37(s6[38],c6[38],andpr9[37],c7[38],s7[37]);


full_add fa7_38(s6[39],c6[39],andpr9[38],c7[39],s7[38]);


full_add fa7_39(s6[40],c6[40],andpr9[39],c7[40],s7[39]);


full_add fa7_40(s6[41],c6[41],andpr9[40],c7[41],s7[40]);


full_add fa7_41(s6[42],c6[42],andpr9[41],c7[42],s7[41]);


full_add fa7_42(s6[43],c6[43],andpr9[42],c7[43],s7[42]);


full_add fa7_43(s6[44],c6[44],andpr9[43],c7[44],s7[43]);


full_add fa7_44(s6[45],c6[45],andpr9[44],c7[45],s7[44]);


full_add fa7_45(s6[46],c6[46],andpr9[45],c7[46],s7[45]);


full_add fa7_46(s6[47],c6[47],andpr9[46],c7[47],s7[46]);


full_add fa7_47(s6[48],c6[48],andpr9[47],c7[48],s7[47]);


full_add fa7_48(s6[49],c6[49],andpr9[48],c7[49],s7[48]);


full_add fa7_49(s6[50],c6[50],andpr9[49],c7[50],s7[49]);


full_add fa7_50(s6[51],c6[51],andpr9[50],c7[51],s7[50]);


full_add fa7_51(s6[52],c6[52],andpr9[51],c7[52],s7[51]);


full_add fa7_52(s6[53],c6[53],andpr9[52],c7[53],s7[52]);


full_add fa7_53(s6[54],c6[54],andpr9[53],c7[54],s7[53]);


full_add fa7_54(s6[55],c6[55],andpr9[54],c7[55],s7[54]);


full_add fa7_55(s6[56],c6[56],andpr9[55],c7[56],s7[55]);


full_add fa7_56(s6[57],c6[57],andpr9[56],c7[57],s7[56]);


full_add fa7_57(s6[58],c6[58],andpr9[57],c7[58],s7[57]);


full_add fa7_58(s6[59],c6[59],andpr9[58],c7[59],s7[58]);


full_add fa7_59(s6[60],c6[60],andpr9[59],c7[60],s7[59]);


full_add fa7_60(s6[61],c6[61],andpr9[60],c7[61],s7[60]);


full_add fa7_61(s6[62],c6[62],andpr9[61],c7[62],s7[61]);


full_add fa7_62(si[7],c6[63],andpr9[62],c7[63],s7[62]);



half_adder ha8(s7[0],c7[0],c8[0],p[8]);


full_add fa8_0(s7[1],c7[1],andpr10[0],c8[1],s8[0]);


full_add fa8_1(s7[2],c7[2],andpr10[1],c8[2],s8[1]);


full_add fa8_2(s7[3],c7[3],andpr10[2],c8[3],s8[2]);


full_add fa8_3(s7[4],c7[4],andpr10[3],c8[4],s8[3]);


full_add fa8_4(s7[5],c7[5],andpr10[4],c8[5],s8[4]);


full_add fa8_5(s7[6],c7[6],andpr10[5],c8[6],s8[5]);


full_add fa8_6(s7[7],c7[7],andpr10[6],c8[7],s8[6]);


full_add fa8_7(s7[8],c7[8],andpr10[7],c8[8],s8[7]);


full_add fa8_8(s7[9],c7[9],andpr10[8],c8[9],s8[8]);


full_add fa8_9(s7[10],c7[10],andpr10[9],c8[10],s8[9]);


full_add fa8_10(s7[11],c7[11],andpr10[10],c8[11],s8[10]);


full_add fa8_11(s7[12],c7[12],andpr10[11],c8[12],s8[11]);


full_add fa8_12(s7[13],c7[13],andpr10[12],c8[13],s8[12]);


full_add fa8_13(s7[14],c7[14],andpr10[13],c8[14],s8[13]);


full_add fa8_14(s7[15],c7[15],andpr10[14],c8[15],s8[14]);


full_add fa8_15(s7[16],c7[16],andpr10[15],c8[16],s8[15]);


full_add fa8_16(s7[17],c7[17],andpr10[16],c8[17],s8[16]);


full_add fa8_17(s7[18],c7[18],andpr10[17],c8[18],s8[17]);


full_add fa8_18(s7[19],c7[19],andpr10[18],c8[19],s8[18]);


full_add fa8_19(s7[20],c7[20],andpr10[19],c8[20],s8[19]);


full_add fa8_20(s7[21],c7[21],andpr10[20],c8[21],s8[20]);


full_add fa8_21(s7[22],c7[22],andpr10[21],c8[22],s8[21]);


full_add fa8_22(s7[23],c7[23],andpr10[22],c8[23],s8[22]);


full_add fa8_23(s7[24],c7[24],andpr10[23],c8[24],s8[23]);


full_add fa8_24(s7[25],c7[25],andpr10[24],c8[25],s8[24]);


full_add fa8_25(s7[26],c7[26],andpr10[25],c8[26],s8[25]);


full_add fa8_26(s7[27],c7[27],andpr10[26],c8[27],s8[26]);


full_add fa8_27(s7[28],c7[28],andpr10[27],c8[28],s8[27]);


full_add fa8_28(s7[29],c7[29],andpr10[28],c8[29],s8[28]);


full_add fa8_29(s7[30],c7[30],andpr10[29],c8[30],s8[29]);


full_add fa8_30(s7[31],c7[31],andpr10[30],c8[31],s8[30]);


full_add fa8_31(s7[32],c7[32],andpr10[31],c8[32],s8[31]);


full_add fa8_32(s7[33],c7[33],andpr10[32],c8[33],s8[32]);


full_add fa8_33(s7[34],c7[34],andpr10[33],c8[34],s8[33]);


full_add fa8_34(s7[35],c7[35],andpr10[34],c8[35],s8[34]);


full_add fa8_35(s7[36],c7[36],andpr10[35],c8[36],s8[35]);


full_add fa8_36(s7[37],c7[37],andpr10[36],c8[37],s8[36]);


full_add fa8_37(s7[38],c7[38],andpr10[37],c8[38],s8[37]);


full_add fa8_38(s7[39],c7[39],andpr10[38],c8[39],s8[38]);


full_add fa8_39(s7[40],c7[40],andpr10[39],c8[40],s8[39]);


full_add fa8_40(s7[41],c7[41],andpr10[40],c8[41],s8[40]);


full_add fa8_41(s7[42],c7[42],andpr10[41],c8[42],s8[41]);


full_add fa8_42(s7[43],c7[43],andpr10[42],c8[43],s8[42]);


full_add fa8_43(s7[44],c7[44],andpr10[43],c8[44],s8[43]);


full_add fa8_44(s7[45],c7[45],andpr10[44],c8[45],s8[44]);


full_add fa8_45(s7[46],c7[46],andpr10[45],c8[46],s8[45]);


full_add fa8_46(s7[47],c7[47],andpr10[46],c8[47],s8[46]);


full_add fa8_47(s7[48],c7[48],andpr10[47],c8[48],s8[47]);


full_add fa8_48(s7[49],c7[49],andpr10[48],c8[49],s8[48]);


full_add fa8_49(s7[50],c7[50],andpr10[49],c8[50],s8[49]);


full_add fa8_50(s7[51],c7[51],andpr10[50],c8[51],s8[50]);


full_add fa8_51(s7[52],c7[52],andpr10[51],c8[52],s8[51]);


full_add fa8_52(s7[53],c7[53],andpr10[52],c8[53],s8[52]);


full_add fa8_53(s7[54],c7[54],andpr10[53],c8[54],s8[53]);


full_add fa8_54(s7[55],c7[55],andpr10[54],c8[55],s8[54]);


full_add fa8_55(s7[56],c7[56],andpr10[55],c8[56],s8[55]);


full_add fa8_56(s7[57],c7[57],andpr10[56],c8[57],s8[56]);


full_add fa8_57(s7[58],c7[58],andpr10[57],c8[58],s8[57]);


full_add fa8_58(s7[59],c7[59],andpr10[58],c8[59],s8[58]);


full_add fa8_59(s7[60],c7[60],andpr10[59],c8[60],s8[59]);


full_add fa8_60(s7[61],c7[61],andpr10[60],c8[61],s8[60]);


full_add fa8_61(s7[62],c7[62],andpr10[61],c8[62],s8[61]);


full_add fa8_62(si[8],c7[63],andpr10[62],c8[63],s8[62]);



half_adder ha9(s8[0],c8[0],c9[0],p[9]);


full_add fa9_0(s8[1],c8[1],andpr11[0],c9[1],s9[0]);


full_add fa9_1(s8[2],c8[2],andpr11[1],c9[2],s9[1]);


full_add fa9_2(s8[3],c8[3],andpr11[2],c9[3],s9[2]);


full_add fa9_3(s8[4],c8[4],andpr11[3],c9[4],s9[3]);


full_add fa9_4(s8[5],c8[5],andpr11[4],c9[5],s9[4]);


full_add fa9_5(s8[6],c8[6],andpr11[5],c9[6],s9[5]);


full_add fa9_6(s8[7],c8[7],andpr11[6],c9[7],s9[6]);


full_add fa9_7(s8[8],c8[8],andpr11[7],c9[8],s9[7]);


full_add fa9_8(s8[9],c8[9],andpr11[8],c9[9],s9[8]);


full_add fa9_9(s8[10],c8[10],andpr11[9],c9[10],s9[9]);


full_add fa9_10(s8[11],c8[11],andpr11[10],c9[11],s9[10]);


full_add fa9_11(s8[12],c8[12],andpr11[11],c9[12],s9[11]);


full_add fa9_12(s8[13],c8[13],andpr11[12],c9[13],s9[12]);


full_add fa9_13(s8[14],c8[14],andpr11[13],c9[14],s9[13]);


full_add fa9_14(s8[15],c8[15],andpr11[14],c9[15],s9[14]);


full_add fa9_15(s8[16],c8[16],andpr11[15],c9[16],s9[15]);


full_add fa9_16(s8[17],c8[17],andpr11[16],c9[17],s9[16]);


full_add fa9_17(s8[18],c8[18],andpr11[17],c9[18],s9[17]);


full_add fa9_18(s8[19],c8[19],andpr11[18],c9[19],s9[18]);


full_add fa9_19(s8[20],c8[20],andpr11[19],c9[20],s9[19]);


full_add fa9_20(s8[21],c8[21],andpr11[20],c9[21],s9[20]);


full_add fa9_21(s8[22],c8[22],andpr11[21],c9[22],s9[21]);


full_add fa9_22(s8[23],c8[23],andpr11[22],c9[23],s9[22]);


full_add fa9_23(s8[24],c8[24],andpr11[23],c9[24],s9[23]);


full_add fa9_24(s8[25],c8[25],andpr11[24],c9[25],s9[24]);


full_add fa9_25(s8[26],c8[26],andpr11[25],c9[26],s9[25]);


full_add fa9_26(s8[27],c8[27],andpr11[26],c9[27],s9[26]);


full_add fa9_27(s8[28],c8[28],andpr11[27],c9[28],s9[27]);


full_add fa9_28(s8[29],c8[29],andpr11[28],c9[29],s9[28]);


full_add fa9_29(s8[30],c8[30],andpr11[29],c9[30],s9[29]);


full_add fa9_30(s8[31],c8[31],andpr11[30],c9[31],s9[30]);


full_add fa9_31(s8[32],c8[32],andpr11[31],c9[32],s9[31]);


full_add fa9_32(s8[33],c8[33],andpr11[32],c9[33],s9[32]);


full_add fa9_33(s8[34],c8[34],andpr11[33],c9[34],s9[33]);


full_add fa9_34(s8[35],c8[35],andpr11[34],c9[35],s9[34]);


full_add fa9_35(s8[36],c8[36],andpr11[35],c9[36],s9[35]);


full_add fa9_36(s8[37],c8[37],andpr11[36],c9[37],s9[36]);


full_add fa9_37(s8[38],c8[38],andpr11[37],c9[38],s9[37]);


full_add fa9_38(s8[39],c8[39],andpr11[38],c9[39],s9[38]);


full_add fa9_39(s8[40],c8[40],andpr11[39],c9[40],s9[39]);


full_add fa9_40(s8[41],c8[41],andpr11[40],c9[41],s9[40]);


full_add fa9_41(s8[42],c8[42],andpr11[41],c9[42],s9[41]);


full_add fa9_42(s8[43],c8[43],andpr11[42],c9[43],s9[42]);


full_add fa9_43(s8[44],c8[44],andpr11[43],c9[44],s9[43]);


full_add fa9_44(s8[45],c8[45],andpr11[44],c9[45],s9[44]);


full_add fa9_45(s8[46],c8[46],andpr11[45],c9[46],s9[45]);


full_add fa9_46(s8[47],c8[47],andpr11[46],c9[47],s9[46]);


full_add fa9_47(s8[48],c8[48],andpr11[47],c9[48],s9[47]);


full_add fa9_48(s8[49],c8[49],andpr11[48],c9[49],s9[48]);


full_add fa9_49(s8[50],c8[50],andpr11[49],c9[50],s9[49]);


full_add fa9_50(s8[51],c8[51],andpr11[50],c9[51],s9[50]);


full_add fa9_51(s8[52],c8[52],andpr11[51],c9[52],s9[51]);


full_add fa9_52(s8[53],c8[53],andpr11[52],c9[53],s9[52]);


full_add fa9_53(s8[54],c8[54],andpr11[53],c9[54],s9[53]);


full_add fa9_54(s8[55],c8[55],andpr11[54],c9[55],s9[54]);


full_add fa9_55(s8[56],c8[56],andpr11[55],c9[56],s9[55]);


full_add fa9_56(s8[57],c8[57],andpr11[56],c9[57],s9[56]);


full_add fa9_57(s8[58],c8[58],andpr11[57],c9[58],s9[57]);


full_add fa9_58(s8[59],c8[59],andpr11[58],c9[59],s9[58]);


full_add fa9_59(s8[60],c8[60],andpr11[59],c9[60],s9[59]);


full_add fa9_60(s8[61],c8[61],andpr11[60],c9[61],s9[60]);


full_add fa9_61(s8[62],c8[62],andpr11[61],c9[62],s9[61]);


full_add fa9_62(si[9],c8[63],andpr11[62],c9[63],s9[62]);



half_adder ha10(s9[0],c9[0],c10[0],p[10]);


full_add fa10_0(s9[1],c9[1],andpr12[0],c10[1],s10[0]);


full_add fa10_1(s9[2],c9[2],andpr12[1],c10[2],s10[1]);


full_add fa10_2(s9[3],c9[3],andpr12[2],c10[3],s10[2]);


full_add fa10_3(s9[4],c9[4],andpr12[3],c10[4],s10[3]);


full_add fa10_4(s9[5],c9[5],andpr12[4],c10[5],s10[4]);


full_add fa10_5(s9[6],c9[6],andpr12[5],c10[6],s10[5]);


full_add fa10_6(s9[7],c9[7],andpr12[6],c10[7],s10[6]);


full_add fa10_7(s9[8],c9[8],andpr12[7],c10[8],s10[7]);


full_add fa10_8(s9[9],c9[9],andpr12[8],c10[9],s10[8]);


full_add fa10_9(s9[10],c9[10],andpr12[9],c10[10],s10[9]);


full_add fa10_10(s9[11],c9[11],andpr12[10],c10[11],s10[10]);


full_add fa10_11(s9[12],c9[12],andpr12[11],c10[12],s10[11]);


full_add fa10_12(s9[13],c9[13],andpr12[12],c10[13],s10[12]);


full_add fa10_13(s9[14],c9[14],andpr12[13],c10[14],s10[13]);


full_add fa10_14(s9[15],c9[15],andpr12[14],c10[15],s10[14]);


full_add fa10_15(s9[16],c9[16],andpr12[15],c10[16],s10[15]);


full_add fa10_16(s9[17],c9[17],andpr12[16],c10[17],s10[16]);


full_add fa10_17(s9[18],c9[18],andpr12[17],c10[18],s10[17]);


full_add fa10_18(s9[19],c9[19],andpr12[18],c10[19],s10[18]);


full_add fa10_19(s9[20],c9[20],andpr12[19],c10[20],s10[19]);


full_add fa10_20(s9[21],c9[21],andpr12[20],c10[21],s10[20]);


full_add fa10_21(s9[22],c9[22],andpr12[21],c10[22],s10[21]);


full_add fa10_22(s9[23],c9[23],andpr12[22],c10[23],s10[22]);


full_add fa10_23(s9[24],c9[24],andpr12[23],c10[24],s10[23]);


full_add fa10_24(s9[25],c9[25],andpr12[24],c10[25],s10[24]);


full_add fa10_25(s9[26],c9[26],andpr12[25],c10[26],s10[25]);


full_add fa10_26(s9[27],c9[27],andpr12[26],c10[27],s10[26]);


full_add fa10_27(s9[28],c9[28],andpr12[27],c10[28],s10[27]);


full_add fa10_28(s9[29],c9[29],andpr12[28],c10[29],s10[28]);


full_add fa10_29(s9[30],c9[30],andpr12[29],c10[30],s10[29]);


full_add fa10_30(s9[31],c9[31],andpr12[30],c10[31],s10[30]);


full_add fa10_31(s9[32],c9[32],andpr12[31],c10[32],s10[31]);


full_add fa10_32(s9[33],c9[33],andpr12[32],c10[33],s10[32]);


full_add fa10_33(s9[34],c9[34],andpr12[33],c10[34],s10[33]);


full_add fa10_34(s9[35],c9[35],andpr12[34],c10[35],s10[34]);


full_add fa10_35(s9[36],c9[36],andpr12[35],c10[36],s10[35]);


full_add fa10_36(s9[37],c9[37],andpr12[36],c10[37],s10[36]);


full_add fa10_37(s9[38],c9[38],andpr12[37],c10[38],s10[37]);


full_add fa10_38(s9[39],c9[39],andpr12[38],c10[39],s10[38]);


full_add fa10_39(s9[40],c9[40],andpr12[39],c10[40],s10[39]);


full_add fa10_40(s9[41],c9[41],andpr12[40],c10[41],s10[40]);


full_add fa10_41(s9[42],c9[42],andpr12[41],c10[42],s10[41]);


full_add fa10_42(s9[43],c9[43],andpr12[42],c10[43],s10[42]);


full_add fa10_43(s9[44],c9[44],andpr12[43],c10[44],s10[43]);


full_add fa10_44(s9[45],c9[45],andpr12[44],c10[45],s10[44]);


full_add fa10_45(s9[46],c9[46],andpr12[45],c10[46],s10[45]);


full_add fa10_46(s9[47],c9[47],andpr12[46],c10[47],s10[46]);


full_add fa10_47(s9[48],c9[48],andpr12[47],c10[48],s10[47]);


full_add fa10_48(s9[49],c9[49],andpr12[48],c10[49],s10[48]);


full_add fa10_49(s9[50],c9[50],andpr12[49],c10[50],s10[49]);


full_add fa10_50(s9[51],c9[51],andpr12[50],c10[51],s10[50]);


full_add fa10_51(s9[52],c9[52],andpr12[51],c10[52],s10[51]);


full_add fa10_52(s9[53],c9[53],andpr12[52],c10[53],s10[52]);


full_add fa10_53(s9[54],c9[54],andpr12[53],c10[54],s10[53]);


full_add fa10_54(s9[55],c9[55],andpr12[54],c10[55],s10[54]);


full_add fa10_55(s9[56],c9[56],andpr12[55],c10[56],s10[55]);


full_add fa10_56(s9[57],c9[57],andpr12[56],c10[57],s10[56]);


full_add fa10_57(s9[58],c9[58],andpr12[57],c10[58],s10[57]);


full_add fa10_58(s9[59],c9[59],andpr12[58],c10[59],s10[58]);


full_add fa10_59(s9[60],c9[60],andpr12[59],c10[60],s10[59]);


full_add fa10_60(s9[61],c9[61],andpr12[60],c10[61],s10[60]);


full_add fa10_61(s9[62],c9[62],andpr12[61],c10[62],s10[61]);


full_add fa10_62(si[10],c9[63],andpr12[62],c10[63],s10[62]);



half_adder ha11(s10[0],c10[0],c11[0],p[11]);


full_add fa11_0(s10[1],c10[1],andpr13[0],c11[1],s11[0]);


full_add fa11_1(s10[2],c10[2],andpr13[1],c11[2],s11[1]);


full_add fa11_2(s10[3],c10[3],andpr13[2],c11[3],s11[2]);


full_add fa11_3(s10[4],c10[4],andpr13[3],c11[4],s11[3]);


full_add fa11_4(s10[5],c10[5],andpr13[4],c11[5],s11[4]);


full_add fa11_5(s10[6],c10[6],andpr13[5],c11[6],s11[5]);


full_add fa11_6(s10[7],c10[7],andpr13[6],c11[7],s11[6]);


full_add fa11_7(s10[8],c10[8],andpr13[7],c11[8],s11[7]);


full_add fa11_8(s10[9],c10[9],andpr13[8],c11[9],s11[8]);


full_add fa11_9(s10[10],c10[10],andpr13[9],c11[10],s11[9]);


full_add fa11_10(s10[11],c10[11],andpr13[10],c11[11],s11[10]);


full_add fa11_11(s10[12],c10[12],andpr13[11],c11[12],s11[11]);


full_add fa11_12(s10[13],c10[13],andpr13[12],c11[13],s11[12]);


full_add fa11_13(s10[14],c10[14],andpr13[13],c11[14],s11[13]);


full_add fa11_14(s10[15],c10[15],andpr13[14],c11[15],s11[14]);


full_add fa11_15(s10[16],c10[16],andpr13[15],c11[16],s11[15]);


full_add fa11_16(s10[17],c10[17],andpr13[16],c11[17],s11[16]);


full_add fa11_17(s10[18],c10[18],andpr13[17],c11[18],s11[17]);


full_add fa11_18(s10[19],c10[19],andpr13[18],c11[19],s11[18]);


full_add fa11_19(s10[20],c10[20],andpr13[19],c11[20],s11[19]);


full_add fa11_20(s10[21],c10[21],andpr13[20],c11[21],s11[20]);


full_add fa11_21(s10[22],c10[22],andpr13[21],c11[22],s11[21]);


full_add fa11_22(s10[23],c10[23],andpr13[22],c11[23],s11[22]);


full_add fa11_23(s10[24],c10[24],andpr13[23],c11[24],s11[23]);


full_add fa11_24(s10[25],c10[25],andpr13[24],c11[25],s11[24]);


full_add fa11_25(s10[26],c10[26],andpr13[25],c11[26],s11[25]);


full_add fa11_26(s10[27],c10[27],andpr13[26],c11[27],s11[26]);


full_add fa11_27(s10[28],c10[28],andpr13[27],c11[28],s11[27]);


full_add fa11_28(s10[29],c10[29],andpr13[28],c11[29],s11[28]);


full_add fa11_29(s10[30],c10[30],andpr13[29],c11[30],s11[29]);


full_add fa11_30(s10[31],c10[31],andpr13[30],c11[31],s11[30]);


full_add fa11_31(s10[32],c10[32],andpr13[31],c11[32],s11[31]);


full_add fa11_32(s10[33],c10[33],andpr13[32],c11[33],s11[32]);


full_add fa11_33(s10[34],c10[34],andpr13[33],c11[34],s11[33]);


full_add fa11_34(s10[35],c10[35],andpr13[34],c11[35],s11[34]);


full_add fa11_35(s10[36],c10[36],andpr13[35],c11[36],s11[35]);


full_add fa11_36(s10[37],c10[37],andpr13[36],c11[37],s11[36]);


full_add fa11_37(s10[38],c10[38],andpr13[37],c11[38],s11[37]);


full_add fa11_38(s10[39],c10[39],andpr13[38],c11[39],s11[38]);


full_add fa11_39(s10[40],c10[40],andpr13[39],c11[40],s11[39]);


full_add fa11_40(s10[41],c10[41],andpr13[40],c11[41],s11[40]);


full_add fa11_41(s10[42],c10[42],andpr13[41],c11[42],s11[41]);


full_add fa11_42(s10[43],c10[43],andpr13[42],c11[43],s11[42]);


full_add fa11_43(s10[44],c10[44],andpr13[43],c11[44],s11[43]);


full_add fa11_44(s10[45],c10[45],andpr13[44],c11[45],s11[44]);


full_add fa11_45(s10[46],c10[46],andpr13[45],c11[46],s11[45]);


full_add fa11_46(s10[47],c10[47],andpr13[46],c11[47],s11[46]);


full_add fa11_47(s10[48],c10[48],andpr13[47],c11[48],s11[47]);


full_add fa11_48(s10[49],c10[49],andpr13[48],c11[49],s11[48]);


full_add fa11_49(s10[50],c10[50],andpr13[49],c11[50],s11[49]);


full_add fa11_50(s10[51],c10[51],andpr13[50],c11[51],s11[50]);


full_add fa11_51(s10[52],c10[52],andpr13[51],c11[52],s11[51]);


full_add fa11_52(s10[53],c10[53],andpr13[52],c11[53],s11[52]);


full_add fa11_53(s10[54],c10[54],andpr13[53],c11[54],s11[53]);


full_add fa11_54(s10[55],c10[55],andpr13[54],c11[55],s11[54]);


full_add fa11_55(s10[56],c10[56],andpr13[55],c11[56],s11[55]);


full_add fa11_56(s10[57],c10[57],andpr13[56],c11[57],s11[56]);


full_add fa11_57(s10[58],c10[58],andpr13[57],c11[58],s11[57]);


full_add fa11_58(s10[59],c10[59],andpr13[58],c11[59],s11[58]);


full_add fa11_59(s10[60],c10[60],andpr13[59],c11[60],s11[59]);


full_add fa11_60(s10[61],c10[61],andpr13[60],c11[61],s11[60]);


full_add fa11_61(s10[62],c10[62],andpr13[61],c11[62],s11[61]);


full_add fa11_62(si[11],c10[63],andpr13[62],c11[63],s11[62]);



half_adder ha12(s11[0],c11[0],c12[0],p[12]);


full_add fa12_0(s11[1],c11[1],andpr14[0],c12[1],s12[0]);


full_add fa12_1(s11[2],c11[2],andpr14[1],c12[2],s12[1]);


full_add fa12_2(s11[3],c11[3],andpr14[2],c12[3],s12[2]);


full_add fa12_3(s11[4],c11[4],andpr14[3],c12[4],s12[3]);


full_add fa12_4(s11[5],c11[5],andpr14[4],c12[5],s12[4]);


full_add fa12_5(s11[6],c11[6],andpr14[5],c12[6],s12[5]);


full_add fa12_6(s11[7],c11[7],andpr14[6],c12[7],s12[6]);


full_add fa12_7(s11[8],c11[8],andpr14[7],c12[8],s12[7]);


full_add fa12_8(s11[9],c11[9],andpr14[8],c12[9],s12[8]);


full_add fa12_9(s11[10],c11[10],andpr14[9],c12[10],s12[9]);


full_add fa12_10(s11[11],c11[11],andpr14[10],c12[11],s12[10]);


full_add fa12_11(s11[12],c11[12],andpr14[11],c12[12],s12[11]);


full_add fa12_12(s11[13],c11[13],andpr14[12],c12[13],s12[12]);


full_add fa12_13(s11[14],c11[14],andpr14[13],c12[14],s12[13]);


full_add fa12_14(s11[15],c11[15],andpr14[14],c12[15],s12[14]);


full_add fa12_15(s11[16],c11[16],andpr14[15],c12[16],s12[15]);


full_add fa12_16(s11[17],c11[17],andpr14[16],c12[17],s12[16]);


full_add fa12_17(s11[18],c11[18],andpr14[17],c12[18],s12[17]);


full_add fa12_18(s11[19],c11[19],andpr14[18],c12[19],s12[18]);


full_add fa12_19(s11[20],c11[20],andpr14[19],c12[20],s12[19]);


full_add fa12_20(s11[21],c11[21],andpr14[20],c12[21],s12[20]);


full_add fa12_21(s11[22],c11[22],andpr14[21],c12[22],s12[21]);


full_add fa12_22(s11[23],c11[23],andpr14[22],c12[23],s12[22]);


full_add fa12_23(s11[24],c11[24],andpr14[23],c12[24],s12[23]);


full_add fa12_24(s11[25],c11[25],andpr14[24],c12[25],s12[24]);


full_add fa12_25(s11[26],c11[26],andpr14[25],c12[26],s12[25]);


full_add fa12_26(s11[27],c11[27],andpr14[26],c12[27],s12[26]);


full_add fa12_27(s11[28],c11[28],andpr14[27],c12[28],s12[27]);


full_add fa12_28(s11[29],c11[29],andpr14[28],c12[29],s12[28]);


full_add fa12_29(s11[30],c11[30],andpr14[29],c12[30],s12[29]);


full_add fa12_30(s11[31],c11[31],andpr14[30],c12[31],s12[30]);


full_add fa12_31(s11[32],c11[32],andpr14[31],c12[32],s12[31]);


full_add fa12_32(s11[33],c11[33],andpr14[32],c12[33],s12[32]);


full_add fa12_33(s11[34],c11[34],andpr14[33],c12[34],s12[33]);


full_add fa12_34(s11[35],c11[35],andpr14[34],c12[35],s12[34]);


full_add fa12_35(s11[36],c11[36],andpr14[35],c12[36],s12[35]);


full_add fa12_36(s11[37],c11[37],andpr14[36],c12[37],s12[36]);


full_add fa12_37(s11[38],c11[38],andpr14[37],c12[38],s12[37]);


full_add fa12_38(s11[39],c11[39],andpr14[38],c12[39],s12[38]);


full_add fa12_39(s11[40],c11[40],andpr14[39],c12[40],s12[39]);


full_add fa12_40(s11[41],c11[41],andpr14[40],c12[41],s12[40]);


full_add fa12_41(s11[42],c11[42],andpr14[41],c12[42],s12[41]);


full_add fa12_42(s11[43],c11[43],andpr14[42],c12[43],s12[42]);


full_add fa12_43(s11[44],c11[44],andpr14[43],c12[44],s12[43]);


full_add fa12_44(s11[45],c11[45],andpr14[44],c12[45],s12[44]);


full_add fa12_45(s11[46],c11[46],andpr14[45],c12[46],s12[45]);


full_add fa12_46(s11[47],c11[47],andpr14[46],c12[47],s12[46]);


full_add fa12_47(s11[48],c11[48],andpr14[47],c12[48],s12[47]);


full_add fa12_48(s11[49],c11[49],andpr14[48],c12[49],s12[48]);


full_add fa12_49(s11[50],c11[50],andpr14[49],c12[50],s12[49]);


full_add fa12_50(s11[51],c11[51],andpr14[50],c12[51],s12[50]);


full_add fa12_51(s11[52],c11[52],andpr14[51],c12[52],s12[51]);


full_add fa12_52(s11[53],c11[53],andpr14[52],c12[53],s12[52]);


full_add fa12_53(s11[54],c11[54],andpr14[53],c12[54],s12[53]);


full_add fa12_54(s11[55],c11[55],andpr14[54],c12[55],s12[54]);


full_add fa12_55(s11[56],c11[56],andpr14[55],c12[56],s12[55]);


full_add fa12_56(s11[57],c11[57],andpr14[56],c12[57],s12[56]);


full_add fa12_57(s11[58],c11[58],andpr14[57],c12[58],s12[57]);


full_add fa12_58(s11[59],c11[59],andpr14[58],c12[59],s12[58]);


full_add fa12_59(s11[60],c11[60],andpr14[59],c12[60],s12[59]);


full_add fa12_60(s11[61],c11[61],andpr14[60],c12[61],s12[60]);


full_add fa12_61(s11[62],c11[62],andpr14[61],c12[62],s12[61]);


full_add fa12_62(si[12],c11[63],andpr14[62],c12[63],s12[62]);



half_adder ha13(s12[0],c12[0],c13[0],p[13]);


full_add fa13_0(s12[1],c12[1],andpr15[0],c13[1],s13[0]);


full_add fa13_1(s12[2],c12[2],andpr15[1],c13[2],s13[1]);


full_add fa13_2(s12[3],c12[3],andpr15[2],c13[3],s13[2]);


full_add fa13_3(s12[4],c12[4],andpr15[3],c13[4],s13[3]);


full_add fa13_4(s12[5],c12[5],andpr15[4],c13[5],s13[4]);


full_add fa13_5(s12[6],c12[6],andpr15[5],c13[6],s13[5]);


full_add fa13_6(s12[7],c12[7],andpr15[6],c13[7],s13[6]);


full_add fa13_7(s12[8],c12[8],andpr15[7],c13[8],s13[7]);


full_add fa13_8(s12[9],c12[9],andpr15[8],c13[9],s13[8]);


full_add fa13_9(s12[10],c12[10],andpr15[9],c13[10],s13[9]);


full_add fa13_10(s12[11],c12[11],andpr15[10],c13[11],s13[10]);


full_add fa13_11(s12[12],c12[12],andpr15[11],c13[12],s13[11]);


full_add fa13_12(s12[13],c12[13],andpr15[12],c13[13],s13[12]);


full_add fa13_13(s12[14],c12[14],andpr15[13],c13[14],s13[13]);


full_add fa13_14(s12[15],c12[15],andpr15[14],c13[15],s13[14]);


full_add fa13_15(s12[16],c12[16],andpr15[15],c13[16],s13[15]);


full_add fa13_16(s12[17],c12[17],andpr15[16],c13[17],s13[16]);


full_add fa13_17(s12[18],c12[18],andpr15[17],c13[18],s13[17]);


full_add fa13_18(s12[19],c12[19],andpr15[18],c13[19],s13[18]);


full_add fa13_19(s12[20],c12[20],andpr15[19],c13[20],s13[19]);


full_add fa13_20(s12[21],c12[21],andpr15[20],c13[21],s13[20]);


full_add fa13_21(s12[22],c12[22],andpr15[21],c13[22],s13[21]);


full_add fa13_22(s12[23],c12[23],andpr15[22],c13[23],s13[22]);


full_add fa13_23(s12[24],c12[24],andpr15[23],c13[24],s13[23]);


full_add fa13_24(s12[25],c12[25],andpr15[24],c13[25],s13[24]);


full_add fa13_25(s12[26],c12[26],andpr15[25],c13[26],s13[25]);


full_add fa13_26(s12[27],c12[27],andpr15[26],c13[27],s13[26]);


full_add fa13_27(s12[28],c12[28],andpr15[27],c13[28],s13[27]);


full_add fa13_28(s12[29],c12[29],andpr15[28],c13[29],s13[28]);


full_add fa13_29(s12[30],c12[30],andpr15[29],c13[30],s13[29]);


full_add fa13_30(s12[31],c12[31],andpr15[30],c13[31],s13[30]);


full_add fa13_31(s12[32],c12[32],andpr15[31],c13[32],s13[31]);


full_add fa13_32(s12[33],c12[33],andpr15[32],c13[33],s13[32]);


full_add fa13_33(s12[34],c12[34],andpr15[33],c13[34],s13[33]);


full_add fa13_34(s12[35],c12[35],andpr15[34],c13[35],s13[34]);


full_add fa13_35(s12[36],c12[36],andpr15[35],c13[36],s13[35]);


full_add fa13_36(s12[37],c12[37],andpr15[36],c13[37],s13[36]);


full_add fa13_37(s12[38],c12[38],andpr15[37],c13[38],s13[37]);


full_add fa13_38(s12[39],c12[39],andpr15[38],c13[39],s13[38]);


full_add fa13_39(s12[40],c12[40],andpr15[39],c13[40],s13[39]);


full_add fa13_40(s12[41],c12[41],andpr15[40],c13[41],s13[40]);


full_add fa13_41(s12[42],c12[42],andpr15[41],c13[42],s13[41]);


full_add fa13_42(s12[43],c12[43],andpr15[42],c13[43],s13[42]);


full_add fa13_43(s12[44],c12[44],andpr15[43],c13[44],s13[43]);


full_add fa13_44(s12[45],c12[45],andpr15[44],c13[45],s13[44]);


full_add fa13_45(s12[46],c12[46],andpr15[45],c13[46],s13[45]);


full_add fa13_46(s12[47],c12[47],andpr15[46],c13[47],s13[46]);


full_add fa13_47(s12[48],c12[48],andpr15[47],c13[48],s13[47]);


full_add fa13_48(s12[49],c12[49],andpr15[48],c13[49],s13[48]);


full_add fa13_49(s12[50],c12[50],andpr15[49],c13[50],s13[49]);


full_add fa13_50(s12[51],c12[51],andpr15[50],c13[51],s13[50]);


full_add fa13_51(s12[52],c12[52],andpr15[51],c13[52],s13[51]);


full_add fa13_52(s12[53],c12[53],andpr15[52],c13[53],s13[52]);


full_add fa13_53(s12[54],c12[54],andpr15[53],c13[54],s13[53]);


full_add fa13_54(s12[55],c12[55],andpr15[54],c13[55],s13[54]);


full_add fa13_55(s12[56],c12[56],andpr15[55],c13[56],s13[55]);


full_add fa13_56(s12[57],c12[57],andpr15[56],c13[57],s13[56]);


full_add fa13_57(s12[58],c12[58],andpr15[57],c13[58],s13[57]);


full_add fa13_58(s12[59],c12[59],andpr15[58],c13[59],s13[58]);


full_add fa13_59(s12[60],c12[60],andpr15[59],c13[60],s13[59]);


full_add fa13_60(s12[61],c12[61],andpr15[60],c13[61],s13[60]);


full_add fa13_61(s12[62],c12[62],andpr15[61],c13[62],s13[61]);


full_add fa13_62(si[13],c12[63],andpr15[62],c13[63],s13[62]);



half_adder ha14(s13[0],c13[0],c14[0],p[14]);


full_add fa14_0(s13[1],c13[1],andpr16[0],c14[1],s14[0]);


full_add fa14_1(s13[2],c13[2],andpr16[1],c14[2],s14[1]);


full_add fa14_2(s13[3],c13[3],andpr16[2],c14[3],s14[2]);


full_add fa14_3(s13[4],c13[4],andpr16[3],c14[4],s14[3]);


full_add fa14_4(s13[5],c13[5],andpr16[4],c14[5],s14[4]);


full_add fa14_5(s13[6],c13[6],andpr16[5],c14[6],s14[5]);


full_add fa14_6(s13[7],c13[7],andpr16[6],c14[7],s14[6]);


full_add fa14_7(s13[8],c13[8],andpr16[7],c14[8],s14[7]);


full_add fa14_8(s13[9],c13[9],andpr16[8],c14[9],s14[8]);


full_add fa14_9(s13[10],c13[10],andpr16[9],c14[10],s14[9]);


full_add fa14_10(s13[11],c13[11],andpr16[10],c14[11],s14[10]);


full_add fa14_11(s13[12],c13[12],andpr16[11],c14[12],s14[11]);


full_add fa14_12(s13[13],c13[13],andpr16[12],c14[13],s14[12]);


full_add fa14_13(s13[14],c13[14],andpr16[13],c14[14],s14[13]);


full_add fa14_14(s13[15],c13[15],andpr16[14],c14[15],s14[14]);


full_add fa14_15(s13[16],c13[16],andpr16[15],c14[16],s14[15]);


full_add fa14_16(s13[17],c13[17],andpr16[16],c14[17],s14[16]);


full_add fa14_17(s13[18],c13[18],andpr16[17],c14[18],s14[17]);


full_add fa14_18(s13[19],c13[19],andpr16[18],c14[19],s14[18]);


full_add fa14_19(s13[20],c13[20],andpr16[19],c14[20],s14[19]);


full_add fa14_20(s13[21],c13[21],andpr16[20],c14[21],s14[20]);


full_add fa14_21(s13[22],c13[22],andpr16[21],c14[22],s14[21]);


full_add fa14_22(s13[23],c13[23],andpr16[22],c14[23],s14[22]);


full_add fa14_23(s13[24],c13[24],andpr16[23],c14[24],s14[23]);


full_add fa14_24(s13[25],c13[25],andpr16[24],c14[25],s14[24]);


full_add fa14_25(s13[26],c13[26],andpr16[25],c14[26],s14[25]);


full_add fa14_26(s13[27],c13[27],andpr16[26],c14[27],s14[26]);


full_add fa14_27(s13[28],c13[28],andpr16[27],c14[28],s14[27]);


full_add fa14_28(s13[29],c13[29],andpr16[28],c14[29],s14[28]);


full_add fa14_29(s13[30],c13[30],andpr16[29],c14[30],s14[29]);


full_add fa14_30(s13[31],c13[31],andpr16[30],c14[31],s14[30]);


full_add fa14_31(s13[32],c13[32],andpr16[31],c14[32],s14[31]);


full_add fa14_32(s13[33],c13[33],andpr16[32],c14[33],s14[32]);


full_add fa14_33(s13[34],c13[34],andpr16[33],c14[34],s14[33]);


full_add fa14_34(s13[35],c13[35],andpr16[34],c14[35],s14[34]);


full_add fa14_35(s13[36],c13[36],andpr16[35],c14[36],s14[35]);


full_add fa14_36(s13[37],c13[37],andpr16[36],c14[37],s14[36]);


full_add fa14_37(s13[38],c13[38],andpr16[37],c14[38],s14[37]);


full_add fa14_38(s13[39],c13[39],andpr16[38],c14[39],s14[38]);


full_add fa14_39(s13[40],c13[40],andpr16[39],c14[40],s14[39]);


full_add fa14_40(s13[41],c13[41],andpr16[40],c14[41],s14[40]);


full_add fa14_41(s13[42],c13[42],andpr16[41],c14[42],s14[41]);


full_add fa14_42(s13[43],c13[43],andpr16[42],c14[43],s14[42]);


full_add fa14_43(s13[44],c13[44],andpr16[43],c14[44],s14[43]);


full_add fa14_44(s13[45],c13[45],andpr16[44],c14[45],s14[44]);


full_add fa14_45(s13[46],c13[46],andpr16[45],c14[46],s14[45]);


full_add fa14_46(s13[47],c13[47],andpr16[46],c14[47],s14[46]);


full_add fa14_47(s13[48],c13[48],andpr16[47],c14[48],s14[47]);


full_add fa14_48(s13[49],c13[49],andpr16[48],c14[49],s14[48]);


full_add fa14_49(s13[50],c13[50],andpr16[49],c14[50],s14[49]);


full_add fa14_50(s13[51],c13[51],andpr16[50],c14[51],s14[50]);


full_add fa14_51(s13[52],c13[52],andpr16[51],c14[52],s14[51]);


full_add fa14_52(s13[53],c13[53],andpr16[52],c14[53],s14[52]);


full_add fa14_53(s13[54],c13[54],andpr16[53],c14[54],s14[53]);


full_add fa14_54(s13[55],c13[55],andpr16[54],c14[55],s14[54]);


full_add fa14_55(s13[56],c13[56],andpr16[55],c14[56],s14[55]);


full_add fa14_56(s13[57],c13[57],andpr16[56],c14[57],s14[56]);


full_add fa14_57(s13[58],c13[58],andpr16[57],c14[58],s14[57]);


full_add fa14_58(s13[59],c13[59],andpr16[58],c14[59],s14[58]);


full_add fa14_59(s13[60],c13[60],andpr16[59],c14[60],s14[59]);


full_add fa14_60(s13[61],c13[61],andpr16[60],c14[61],s14[60]);


full_add fa14_61(s13[62],c13[62],andpr16[61],c14[62],s14[61]);


full_add fa14_62(si[14],c13[63],andpr16[62],c14[63],s14[62]);



half_adder ha15(s14[0],c14[0],c15[0],p[15]);


full_add fa15_0(s14[1],c14[1],andpr17[0],c15[1],s15[0]);


full_add fa15_1(s14[2],c14[2],andpr17[1],c15[2],s15[1]);


full_add fa15_2(s14[3],c14[3],andpr17[2],c15[3],s15[2]);


full_add fa15_3(s14[4],c14[4],andpr17[3],c15[4],s15[3]);


full_add fa15_4(s14[5],c14[5],andpr17[4],c15[5],s15[4]);


full_add fa15_5(s14[6],c14[6],andpr17[5],c15[6],s15[5]);


full_add fa15_6(s14[7],c14[7],andpr17[6],c15[7],s15[6]);


full_add fa15_7(s14[8],c14[8],andpr17[7],c15[8],s15[7]);


full_add fa15_8(s14[9],c14[9],andpr17[8],c15[9],s15[8]);


full_add fa15_9(s14[10],c14[10],andpr17[9],c15[10],s15[9]);


full_add fa15_10(s14[11],c14[11],andpr17[10],c15[11],s15[10]);


full_add fa15_11(s14[12],c14[12],andpr17[11],c15[12],s15[11]);


full_add fa15_12(s14[13],c14[13],andpr17[12],c15[13],s15[12]);


full_add fa15_13(s14[14],c14[14],andpr17[13],c15[14],s15[13]);


full_add fa15_14(s14[15],c14[15],andpr17[14],c15[15],s15[14]);


full_add fa15_15(s14[16],c14[16],andpr17[15],c15[16],s15[15]);


full_add fa15_16(s14[17],c14[17],andpr17[16],c15[17],s15[16]);


full_add fa15_17(s14[18],c14[18],andpr17[17],c15[18],s15[17]);


full_add fa15_18(s14[19],c14[19],andpr17[18],c15[19],s15[18]);


full_add fa15_19(s14[20],c14[20],andpr17[19],c15[20],s15[19]);


full_add fa15_20(s14[21],c14[21],andpr17[20],c15[21],s15[20]);


full_add fa15_21(s14[22],c14[22],andpr17[21],c15[22],s15[21]);


full_add fa15_22(s14[23],c14[23],andpr17[22],c15[23],s15[22]);


full_add fa15_23(s14[24],c14[24],andpr17[23],c15[24],s15[23]);


full_add fa15_24(s14[25],c14[25],andpr17[24],c15[25],s15[24]);


full_add fa15_25(s14[26],c14[26],andpr17[25],c15[26],s15[25]);


full_add fa15_26(s14[27],c14[27],andpr17[26],c15[27],s15[26]);


full_add fa15_27(s14[28],c14[28],andpr17[27],c15[28],s15[27]);


full_add fa15_28(s14[29],c14[29],andpr17[28],c15[29],s15[28]);


full_add fa15_29(s14[30],c14[30],andpr17[29],c15[30],s15[29]);


full_add fa15_30(s14[31],c14[31],andpr17[30],c15[31],s15[30]);


full_add fa15_31(s14[32],c14[32],andpr17[31],c15[32],s15[31]);


full_add fa15_32(s14[33],c14[33],andpr17[32],c15[33],s15[32]);


full_add fa15_33(s14[34],c14[34],andpr17[33],c15[34],s15[33]);


full_add fa15_34(s14[35],c14[35],andpr17[34],c15[35],s15[34]);


full_add fa15_35(s14[36],c14[36],andpr17[35],c15[36],s15[35]);


full_add fa15_36(s14[37],c14[37],andpr17[36],c15[37],s15[36]);


full_add fa15_37(s14[38],c14[38],andpr17[37],c15[38],s15[37]);


full_add fa15_38(s14[39],c14[39],andpr17[38],c15[39],s15[38]);


full_add fa15_39(s14[40],c14[40],andpr17[39],c15[40],s15[39]);


full_add fa15_40(s14[41],c14[41],andpr17[40],c15[41],s15[40]);


full_add fa15_41(s14[42],c14[42],andpr17[41],c15[42],s15[41]);


full_add fa15_42(s14[43],c14[43],andpr17[42],c15[43],s15[42]);


full_add fa15_43(s14[44],c14[44],andpr17[43],c15[44],s15[43]);


full_add fa15_44(s14[45],c14[45],andpr17[44],c15[45],s15[44]);


full_add fa15_45(s14[46],c14[46],andpr17[45],c15[46],s15[45]);


full_add fa15_46(s14[47],c14[47],andpr17[46],c15[47],s15[46]);


full_add fa15_47(s14[48],c14[48],andpr17[47],c15[48],s15[47]);


full_add fa15_48(s14[49],c14[49],andpr17[48],c15[49],s15[48]);


full_add fa15_49(s14[50],c14[50],andpr17[49],c15[50],s15[49]);


full_add fa15_50(s14[51],c14[51],andpr17[50],c15[51],s15[50]);


full_add fa15_51(s14[52],c14[52],andpr17[51],c15[52],s15[51]);


full_add fa15_52(s14[53],c14[53],andpr17[52],c15[53],s15[52]);


full_add fa15_53(s14[54],c14[54],andpr17[53],c15[54],s15[53]);


full_add fa15_54(s14[55],c14[55],andpr17[54],c15[55],s15[54]);


full_add fa15_55(s14[56],c14[56],andpr17[55],c15[56],s15[55]);


full_add fa15_56(s14[57],c14[57],andpr17[56],c15[57],s15[56]);


full_add fa15_57(s14[58],c14[58],andpr17[57],c15[58],s15[57]);


full_add fa15_58(s14[59],c14[59],andpr17[58],c15[59],s15[58]);


full_add fa15_59(s14[60],c14[60],andpr17[59],c15[60],s15[59]);


full_add fa15_60(s14[61],c14[61],andpr17[60],c15[61],s15[60]);


full_add fa15_61(s14[62],c14[62],andpr17[61],c15[62],s15[61]);


full_add fa15_62(si[15],c14[63],andpr17[62],c15[63],s15[62]);



half_adder ha16(s15[0],c15[0],c16[0],p[16]);


full_add fa16_0(s15[1],c15[1],andpr18[0],c16[1],s16[0]);


full_add fa16_1(s15[2],c15[2],andpr18[1],c16[2],s16[1]);


full_add fa16_2(s15[3],c15[3],andpr18[2],c16[3],s16[2]);


full_add fa16_3(s15[4],c15[4],andpr18[3],c16[4],s16[3]);


full_add fa16_4(s15[5],c15[5],andpr18[4],c16[5],s16[4]);


full_add fa16_5(s15[6],c15[6],andpr18[5],c16[6],s16[5]);


full_add fa16_6(s15[7],c15[7],andpr18[6],c16[7],s16[6]);


full_add fa16_7(s15[8],c15[8],andpr18[7],c16[8],s16[7]);


full_add fa16_8(s15[9],c15[9],andpr18[8],c16[9],s16[8]);


full_add fa16_9(s15[10],c15[10],andpr18[9],c16[10],s16[9]);


full_add fa16_10(s15[11],c15[11],andpr18[10],c16[11],s16[10]);


full_add fa16_11(s15[12],c15[12],andpr18[11],c16[12],s16[11]);


full_add fa16_12(s15[13],c15[13],andpr18[12],c16[13],s16[12]);


full_add fa16_13(s15[14],c15[14],andpr18[13],c16[14],s16[13]);


full_add fa16_14(s15[15],c15[15],andpr18[14],c16[15],s16[14]);


full_add fa16_15(s15[16],c15[16],andpr18[15],c16[16],s16[15]);


full_add fa16_16(s15[17],c15[17],andpr18[16],c16[17],s16[16]);


full_add fa16_17(s15[18],c15[18],andpr18[17],c16[18],s16[17]);


full_add fa16_18(s15[19],c15[19],andpr18[18],c16[19],s16[18]);


full_add fa16_19(s15[20],c15[20],andpr18[19],c16[20],s16[19]);


full_add fa16_20(s15[21],c15[21],andpr18[20],c16[21],s16[20]);


full_add fa16_21(s15[22],c15[22],andpr18[21],c16[22],s16[21]);


full_add fa16_22(s15[23],c15[23],andpr18[22],c16[23],s16[22]);


full_add fa16_23(s15[24],c15[24],andpr18[23],c16[24],s16[23]);


full_add fa16_24(s15[25],c15[25],andpr18[24],c16[25],s16[24]);


full_add fa16_25(s15[26],c15[26],andpr18[25],c16[26],s16[25]);


full_add fa16_26(s15[27],c15[27],andpr18[26],c16[27],s16[26]);


full_add fa16_27(s15[28],c15[28],andpr18[27],c16[28],s16[27]);


full_add fa16_28(s15[29],c15[29],andpr18[28],c16[29],s16[28]);


full_add fa16_29(s15[30],c15[30],andpr18[29],c16[30],s16[29]);


full_add fa16_30(s15[31],c15[31],andpr18[30],c16[31],s16[30]);


full_add fa16_31(s15[32],c15[32],andpr18[31],c16[32],s16[31]);


full_add fa16_32(s15[33],c15[33],andpr18[32],c16[33],s16[32]);


full_add fa16_33(s15[34],c15[34],andpr18[33],c16[34],s16[33]);


full_add fa16_34(s15[35],c15[35],andpr18[34],c16[35],s16[34]);


full_add fa16_35(s15[36],c15[36],andpr18[35],c16[36],s16[35]);


full_add fa16_36(s15[37],c15[37],andpr18[36],c16[37],s16[36]);


full_add fa16_37(s15[38],c15[38],andpr18[37],c16[38],s16[37]);


full_add fa16_38(s15[39],c15[39],andpr18[38],c16[39],s16[38]);


full_add fa16_39(s15[40],c15[40],andpr18[39],c16[40],s16[39]);


full_add fa16_40(s15[41],c15[41],andpr18[40],c16[41],s16[40]);


full_add fa16_41(s15[42],c15[42],andpr18[41],c16[42],s16[41]);


full_add fa16_42(s15[43],c15[43],andpr18[42],c16[43],s16[42]);


full_add fa16_43(s15[44],c15[44],andpr18[43],c16[44],s16[43]);


full_add fa16_44(s15[45],c15[45],andpr18[44],c16[45],s16[44]);


full_add fa16_45(s15[46],c15[46],andpr18[45],c16[46],s16[45]);


full_add fa16_46(s15[47],c15[47],andpr18[46],c16[47],s16[46]);


full_add fa16_47(s15[48],c15[48],andpr18[47],c16[48],s16[47]);


full_add fa16_48(s15[49],c15[49],andpr18[48],c16[49],s16[48]);


full_add fa16_49(s15[50],c15[50],andpr18[49],c16[50],s16[49]);


full_add fa16_50(s15[51],c15[51],andpr18[50],c16[51],s16[50]);


full_add fa16_51(s15[52],c15[52],andpr18[51],c16[52],s16[51]);


full_add fa16_52(s15[53],c15[53],andpr18[52],c16[53],s16[52]);


full_add fa16_53(s15[54],c15[54],andpr18[53],c16[54],s16[53]);


full_add fa16_54(s15[55],c15[55],andpr18[54],c16[55],s16[54]);


full_add fa16_55(s15[56],c15[56],andpr18[55],c16[56],s16[55]);


full_add fa16_56(s15[57],c15[57],andpr18[56],c16[57],s16[56]);


full_add fa16_57(s15[58],c15[58],andpr18[57],c16[58],s16[57]);


full_add fa16_58(s15[59],c15[59],andpr18[58],c16[59],s16[58]);


full_add fa16_59(s15[60],c15[60],andpr18[59],c16[60],s16[59]);


full_add fa16_60(s15[61],c15[61],andpr18[60],c16[61],s16[60]);


full_add fa16_61(s15[62],c15[62],andpr18[61],c16[62],s16[61]);


full_add fa16_62(si[16],c15[63],andpr18[62],c16[63],s16[62]);



half_adder ha17(s16[0],c16[0],c17[0],p[17]);


full_add fa17_0(s16[1],c16[1],andpr19[0],c17[1],s17[0]);


full_add fa17_1(s16[2],c16[2],andpr19[1],c17[2],s17[1]);


full_add fa17_2(s16[3],c16[3],andpr19[2],c17[3],s17[2]);


full_add fa17_3(s16[4],c16[4],andpr19[3],c17[4],s17[3]);


full_add fa17_4(s16[5],c16[5],andpr19[4],c17[5],s17[4]);


full_add fa17_5(s16[6],c16[6],andpr19[5],c17[6],s17[5]);


full_add fa17_6(s16[7],c16[7],andpr19[6],c17[7],s17[6]);


full_add fa17_7(s16[8],c16[8],andpr19[7],c17[8],s17[7]);


full_add fa17_8(s16[9],c16[9],andpr19[8],c17[9],s17[8]);


full_add fa17_9(s16[10],c16[10],andpr19[9],c17[10],s17[9]);


full_add fa17_10(s16[11],c16[11],andpr19[10],c17[11],s17[10]);


full_add fa17_11(s16[12],c16[12],andpr19[11],c17[12],s17[11]);


full_add fa17_12(s16[13],c16[13],andpr19[12],c17[13],s17[12]);


full_add fa17_13(s16[14],c16[14],andpr19[13],c17[14],s17[13]);


full_add fa17_14(s16[15],c16[15],andpr19[14],c17[15],s17[14]);


full_add fa17_15(s16[16],c16[16],andpr19[15],c17[16],s17[15]);


full_add fa17_16(s16[17],c16[17],andpr19[16],c17[17],s17[16]);


full_add fa17_17(s16[18],c16[18],andpr19[17],c17[18],s17[17]);


full_add fa17_18(s16[19],c16[19],andpr19[18],c17[19],s17[18]);


full_add fa17_19(s16[20],c16[20],andpr19[19],c17[20],s17[19]);


full_add fa17_20(s16[21],c16[21],andpr19[20],c17[21],s17[20]);


full_add fa17_21(s16[22],c16[22],andpr19[21],c17[22],s17[21]);


full_add fa17_22(s16[23],c16[23],andpr19[22],c17[23],s17[22]);


full_add fa17_23(s16[24],c16[24],andpr19[23],c17[24],s17[23]);


full_add fa17_24(s16[25],c16[25],andpr19[24],c17[25],s17[24]);


full_add fa17_25(s16[26],c16[26],andpr19[25],c17[26],s17[25]);


full_add fa17_26(s16[27],c16[27],andpr19[26],c17[27],s17[26]);


full_add fa17_27(s16[28],c16[28],andpr19[27],c17[28],s17[27]);


full_add fa17_28(s16[29],c16[29],andpr19[28],c17[29],s17[28]);


full_add fa17_29(s16[30],c16[30],andpr19[29],c17[30],s17[29]);


full_add fa17_30(s16[31],c16[31],andpr19[30],c17[31],s17[30]);


full_add fa17_31(s16[32],c16[32],andpr19[31],c17[32],s17[31]);


full_add fa17_32(s16[33],c16[33],andpr19[32],c17[33],s17[32]);


full_add fa17_33(s16[34],c16[34],andpr19[33],c17[34],s17[33]);


full_add fa17_34(s16[35],c16[35],andpr19[34],c17[35],s17[34]);


full_add fa17_35(s16[36],c16[36],andpr19[35],c17[36],s17[35]);


full_add fa17_36(s16[37],c16[37],andpr19[36],c17[37],s17[36]);


full_add fa17_37(s16[38],c16[38],andpr19[37],c17[38],s17[37]);


full_add fa17_38(s16[39],c16[39],andpr19[38],c17[39],s17[38]);


full_add fa17_39(s16[40],c16[40],andpr19[39],c17[40],s17[39]);


full_add fa17_40(s16[41],c16[41],andpr19[40],c17[41],s17[40]);


full_add fa17_41(s16[42],c16[42],andpr19[41],c17[42],s17[41]);


full_add fa17_42(s16[43],c16[43],andpr19[42],c17[43],s17[42]);


full_add fa17_43(s16[44],c16[44],andpr19[43],c17[44],s17[43]);


full_add fa17_44(s16[45],c16[45],andpr19[44],c17[45],s17[44]);


full_add fa17_45(s16[46],c16[46],andpr19[45],c17[46],s17[45]);


full_add fa17_46(s16[47],c16[47],andpr19[46],c17[47],s17[46]);


full_add fa17_47(s16[48],c16[48],andpr19[47],c17[48],s17[47]);


full_add fa17_48(s16[49],c16[49],andpr19[48],c17[49],s17[48]);


full_add fa17_49(s16[50],c16[50],andpr19[49],c17[50],s17[49]);


full_add fa17_50(s16[51],c16[51],andpr19[50],c17[51],s17[50]);


full_add fa17_51(s16[52],c16[52],andpr19[51],c17[52],s17[51]);


full_add fa17_52(s16[53],c16[53],andpr19[52],c17[53],s17[52]);


full_add fa17_53(s16[54],c16[54],andpr19[53],c17[54],s17[53]);


full_add fa17_54(s16[55],c16[55],andpr19[54],c17[55],s17[54]);


full_add fa17_55(s16[56],c16[56],andpr19[55],c17[56],s17[55]);


full_add fa17_56(s16[57],c16[57],andpr19[56],c17[57],s17[56]);


full_add fa17_57(s16[58],c16[58],andpr19[57],c17[58],s17[57]);


full_add fa17_58(s16[59],c16[59],andpr19[58],c17[59],s17[58]);


full_add fa17_59(s16[60],c16[60],andpr19[59],c17[60],s17[59]);


full_add fa17_60(s16[61],c16[61],andpr19[60],c17[61],s17[60]);


full_add fa17_61(s16[62],c16[62],andpr19[61],c17[62],s17[61]);


full_add fa17_62(si[17],c16[63],andpr19[62],c17[63],s17[62]);



half_adder ha18(s17[0],c17[0],c18[0],p[18]);


full_add fa18_0(s17[1],c17[1],andpr20[0],c18[1],s18[0]);


full_add fa18_1(s17[2],c17[2],andpr20[1],c18[2],s18[1]);


full_add fa18_2(s17[3],c17[3],andpr20[2],c18[3],s18[2]);


full_add fa18_3(s17[4],c17[4],andpr20[3],c18[4],s18[3]);


full_add fa18_4(s17[5],c17[5],andpr20[4],c18[5],s18[4]);


full_add fa18_5(s17[6],c17[6],andpr20[5],c18[6],s18[5]);


full_add fa18_6(s17[7],c17[7],andpr20[6],c18[7],s18[6]);


full_add fa18_7(s17[8],c17[8],andpr20[7],c18[8],s18[7]);


full_add fa18_8(s17[9],c17[9],andpr20[8],c18[9],s18[8]);


full_add fa18_9(s17[10],c17[10],andpr20[9],c18[10],s18[9]);


full_add fa18_10(s17[11],c17[11],andpr20[10],c18[11],s18[10]);


full_add fa18_11(s17[12],c17[12],andpr20[11],c18[12],s18[11]);


full_add fa18_12(s17[13],c17[13],andpr20[12],c18[13],s18[12]);


full_add fa18_13(s17[14],c17[14],andpr20[13],c18[14],s18[13]);


full_add fa18_14(s17[15],c17[15],andpr20[14],c18[15],s18[14]);


full_add fa18_15(s17[16],c17[16],andpr20[15],c18[16],s18[15]);


full_add fa18_16(s17[17],c17[17],andpr20[16],c18[17],s18[16]);


full_add fa18_17(s17[18],c17[18],andpr20[17],c18[18],s18[17]);


full_add fa18_18(s17[19],c17[19],andpr20[18],c18[19],s18[18]);


full_add fa18_19(s17[20],c17[20],andpr20[19],c18[20],s18[19]);


full_add fa18_20(s17[21],c17[21],andpr20[20],c18[21],s18[20]);


full_add fa18_21(s17[22],c17[22],andpr20[21],c18[22],s18[21]);


full_add fa18_22(s17[23],c17[23],andpr20[22],c18[23],s18[22]);


full_add fa18_23(s17[24],c17[24],andpr20[23],c18[24],s18[23]);


full_add fa18_24(s17[25],c17[25],andpr20[24],c18[25],s18[24]);


full_add fa18_25(s17[26],c17[26],andpr20[25],c18[26],s18[25]);


full_add fa18_26(s17[27],c17[27],andpr20[26],c18[27],s18[26]);


full_add fa18_27(s17[28],c17[28],andpr20[27],c18[28],s18[27]);


full_add fa18_28(s17[29],c17[29],andpr20[28],c18[29],s18[28]);


full_add fa18_29(s17[30],c17[30],andpr20[29],c18[30],s18[29]);


full_add fa18_30(s17[31],c17[31],andpr20[30],c18[31],s18[30]);


full_add fa18_31(s17[32],c17[32],andpr20[31],c18[32],s18[31]);


full_add fa18_32(s17[33],c17[33],andpr20[32],c18[33],s18[32]);


full_add fa18_33(s17[34],c17[34],andpr20[33],c18[34],s18[33]);


full_add fa18_34(s17[35],c17[35],andpr20[34],c18[35],s18[34]);


full_add fa18_35(s17[36],c17[36],andpr20[35],c18[36],s18[35]);


full_add fa18_36(s17[37],c17[37],andpr20[36],c18[37],s18[36]);


full_add fa18_37(s17[38],c17[38],andpr20[37],c18[38],s18[37]);


full_add fa18_38(s17[39],c17[39],andpr20[38],c18[39],s18[38]);


full_add fa18_39(s17[40],c17[40],andpr20[39],c18[40],s18[39]);


full_add fa18_40(s17[41],c17[41],andpr20[40],c18[41],s18[40]);


full_add fa18_41(s17[42],c17[42],andpr20[41],c18[42],s18[41]);


full_add fa18_42(s17[43],c17[43],andpr20[42],c18[43],s18[42]);


full_add fa18_43(s17[44],c17[44],andpr20[43],c18[44],s18[43]);


full_add fa18_44(s17[45],c17[45],andpr20[44],c18[45],s18[44]);


full_add fa18_45(s17[46],c17[46],andpr20[45],c18[46],s18[45]);


full_add fa18_46(s17[47],c17[47],andpr20[46],c18[47],s18[46]);


full_add fa18_47(s17[48],c17[48],andpr20[47],c18[48],s18[47]);


full_add fa18_48(s17[49],c17[49],andpr20[48],c18[49],s18[48]);


full_add fa18_49(s17[50],c17[50],andpr20[49],c18[50],s18[49]);


full_add fa18_50(s17[51],c17[51],andpr20[50],c18[51],s18[50]);


full_add fa18_51(s17[52],c17[52],andpr20[51],c18[52],s18[51]);


full_add fa18_52(s17[53],c17[53],andpr20[52],c18[53],s18[52]);


full_add fa18_53(s17[54],c17[54],andpr20[53],c18[54],s18[53]);


full_add fa18_54(s17[55],c17[55],andpr20[54],c18[55],s18[54]);


full_add fa18_55(s17[56],c17[56],andpr20[55],c18[56],s18[55]);


full_add fa18_56(s17[57],c17[57],andpr20[56],c18[57],s18[56]);


full_add fa18_57(s17[58],c17[58],andpr20[57],c18[58],s18[57]);


full_add fa18_58(s17[59],c17[59],andpr20[58],c18[59],s18[58]);


full_add fa18_59(s17[60],c17[60],andpr20[59],c18[60],s18[59]);


full_add fa18_60(s17[61],c17[61],andpr20[60],c18[61],s18[60]);


full_add fa18_61(s17[62],c17[62],andpr20[61],c18[62],s18[61]);


full_add fa18_62(si[18],c17[63],andpr20[62],c18[63],s18[62]);



half_adder ha19(s18[0],c18[0],c19[0],p[19]);


full_add fa19_0(s18[1],c18[1],andpr21[0],c19[1],s19[0]);


full_add fa19_1(s18[2],c18[2],andpr21[1],c19[2],s19[1]);


full_add fa19_2(s18[3],c18[3],andpr21[2],c19[3],s19[2]);


full_add fa19_3(s18[4],c18[4],andpr21[3],c19[4],s19[3]);


full_add fa19_4(s18[5],c18[5],andpr21[4],c19[5],s19[4]);


full_add fa19_5(s18[6],c18[6],andpr21[5],c19[6],s19[5]);


full_add fa19_6(s18[7],c18[7],andpr21[6],c19[7],s19[6]);


full_add fa19_7(s18[8],c18[8],andpr21[7],c19[8],s19[7]);


full_add fa19_8(s18[9],c18[9],andpr21[8],c19[9],s19[8]);


full_add fa19_9(s18[10],c18[10],andpr21[9],c19[10],s19[9]);


full_add fa19_10(s18[11],c18[11],andpr21[10],c19[11],s19[10]);


full_add fa19_11(s18[12],c18[12],andpr21[11],c19[12],s19[11]);


full_add fa19_12(s18[13],c18[13],andpr21[12],c19[13],s19[12]);


full_add fa19_13(s18[14],c18[14],andpr21[13],c19[14],s19[13]);


full_add fa19_14(s18[15],c18[15],andpr21[14],c19[15],s19[14]);


full_add fa19_15(s18[16],c18[16],andpr21[15],c19[16],s19[15]);


full_add fa19_16(s18[17],c18[17],andpr21[16],c19[17],s19[16]);


full_add fa19_17(s18[18],c18[18],andpr21[17],c19[18],s19[17]);


full_add fa19_18(s18[19],c18[19],andpr21[18],c19[19],s19[18]);


full_add fa19_19(s18[20],c18[20],andpr21[19],c19[20],s19[19]);


full_add fa19_20(s18[21],c18[21],andpr21[20],c19[21],s19[20]);


full_add fa19_21(s18[22],c18[22],andpr21[21],c19[22],s19[21]);


full_add fa19_22(s18[23],c18[23],andpr21[22],c19[23],s19[22]);


full_add fa19_23(s18[24],c18[24],andpr21[23],c19[24],s19[23]);


full_add fa19_24(s18[25],c18[25],andpr21[24],c19[25],s19[24]);


full_add fa19_25(s18[26],c18[26],andpr21[25],c19[26],s19[25]);


full_add fa19_26(s18[27],c18[27],andpr21[26],c19[27],s19[26]);


full_add fa19_27(s18[28],c18[28],andpr21[27],c19[28],s19[27]);


full_add fa19_28(s18[29],c18[29],andpr21[28],c19[29],s19[28]);


full_add fa19_29(s18[30],c18[30],andpr21[29],c19[30],s19[29]);


full_add fa19_30(s18[31],c18[31],andpr21[30],c19[31],s19[30]);


full_add fa19_31(s18[32],c18[32],andpr21[31],c19[32],s19[31]);


full_add fa19_32(s18[33],c18[33],andpr21[32],c19[33],s19[32]);


full_add fa19_33(s18[34],c18[34],andpr21[33],c19[34],s19[33]);


full_add fa19_34(s18[35],c18[35],andpr21[34],c19[35],s19[34]);


full_add fa19_35(s18[36],c18[36],andpr21[35],c19[36],s19[35]);


full_add fa19_36(s18[37],c18[37],andpr21[36],c19[37],s19[36]);


full_add fa19_37(s18[38],c18[38],andpr21[37],c19[38],s19[37]);


full_add fa19_38(s18[39],c18[39],andpr21[38],c19[39],s19[38]);


full_add fa19_39(s18[40],c18[40],andpr21[39],c19[40],s19[39]);


full_add fa19_40(s18[41],c18[41],andpr21[40],c19[41],s19[40]);


full_add fa19_41(s18[42],c18[42],andpr21[41],c19[42],s19[41]);


full_add fa19_42(s18[43],c18[43],andpr21[42],c19[43],s19[42]);


full_add fa19_43(s18[44],c18[44],andpr21[43],c19[44],s19[43]);


full_add fa19_44(s18[45],c18[45],andpr21[44],c19[45],s19[44]);


full_add fa19_45(s18[46],c18[46],andpr21[45],c19[46],s19[45]);


full_add fa19_46(s18[47],c18[47],andpr21[46],c19[47],s19[46]);


full_add fa19_47(s18[48],c18[48],andpr21[47],c19[48],s19[47]);


full_add fa19_48(s18[49],c18[49],andpr21[48],c19[49],s19[48]);


full_add fa19_49(s18[50],c18[50],andpr21[49],c19[50],s19[49]);


full_add fa19_50(s18[51],c18[51],andpr21[50],c19[51],s19[50]);


full_add fa19_51(s18[52],c18[52],andpr21[51],c19[52],s19[51]);


full_add fa19_52(s18[53],c18[53],andpr21[52],c19[53],s19[52]);


full_add fa19_53(s18[54],c18[54],andpr21[53],c19[54],s19[53]);


full_add fa19_54(s18[55],c18[55],andpr21[54],c19[55],s19[54]);


full_add fa19_55(s18[56],c18[56],andpr21[55],c19[56],s19[55]);


full_add fa19_56(s18[57],c18[57],andpr21[56],c19[57],s19[56]);


full_add fa19_57(s18[58],c18[58],andpr21[57],c19[58],s19[57]);


full_add fa19_58(s18[59],c18[59],andpr21[58],c19[59],s19[58]);


full_add fa19_59(s18[60],c18[60],andpr21[59],c19[60],s19[59]);


full_add fa19_60(s18[61],c18[61],andpr21[60],c19[61],s19[60]);


full_add fa19_61(s18[62],c18[62],andpr21[61],c19[62],s19[61]);


full_add fa19_62(si[19],c18[63],andpr21[62],c19[63],s19[62]);



half_adder ha20(s19[0],c19[0],c20[0],p[20]);


full_add fa20_0(s19[1],c19[1],andpr22[0],c20[1],s20[0]);


full_add fa20_1(s19[2],c19[2],andpr22[1],c20[2],s20[1]);


full_add fa20_2(s19[3],c19[3],andpr22[2],c20[3],s20[2]);


full_add fa20_3(s19[4],c19[4],andpr22[3],c20[4],s20[3]);


full_add fa20_4(s19[5],c19[5],andpr22[4],c20[5],s20[4]);


full_add fa20_5(s19[6],c19[6],andpr22[5],c20[6],s20[5]);


full_add fa20_6(s19[7],c19[7],andpr22[6],c20[7],s20[6]);


full_add fa20_7(s19[8],c19[8],andpr22[7],c20[8],s20[7]);


full_add fa20_8(s19[9],c19[9],andpr22[8],c20[9],s20[8]);


full_add fa20_9(s19[10],c19[10],andpr22[9],c20[10],s20[9]);


full_add fa20_10(s19[11],c19[11],andpr22[10],c20[11],s20[10]);


full_add fa20_11(s19[12],c19[12],andpr22[11],c20[12],s20[11]);


full_add fa20_12(s19[13],c19[13],andpr22[12],c20[13],s20[12]);


full_add fa20_13(s19[14],c19[14],andpr22[13],c20[14],s20[13]);


full_add fa20_14(s19[15],c19[15],andpr22[14],c20[15],s20[14]);


full_add fa20_15(s19[16],c19[16],andpr22[15],c20[16],s20[15]);


full_add fa20_16(s19[17],c19[17],andpr22[16],c20[17],s20[16]);


full_add fa20_17(s19[18],c19[18],andpr22[17],c20[18],s20[17]);


full_add fa20_18(s19[19],c19[19],andpr22[18],c20[19],s20[18]);


full_add fa20_19(s19[20],c19[20],andpr22[19],c20[20],s20[19]);


full_add fa20_20(s19[21],c19[21],andpr22[20],c20[21],s20[20]);


full_add fa20_21(s19[22],c19[22],andpr22[21],c20[22],s20[21]);


full_add fa20_22(s19[23],c19[23],andpr22[22],c20[23],s20[22]);


full_add fa20_23(s19[24],c19[24],andpr22[23],c20[24],s20[23]);


full_add fa20_24(s19[25],c19[25],andpr22[24],c20[25],s20[24]);


full_add fa20_25(s19[26],c19[26],andpr22[25],c20[26],s20[25]);


full_add fa20_26(s19[27],c19[27],andpr22[26],c20[27],s20[26]);


full_add fa20_27(s19[28],c19[28],andpr22[27],c20[28],s20[27]);


full_add fa20_28(s19[29],c19[29],andpr22[28],c20[29],s20[28]);


full_add fa20_29(s19[30],c19[30],andpr22[29],c20[30],s20[29]);


full_add fa20_30(s19[31],c19[31],andpr22[30],c20[31],s20[30]);


full_add fa20_31(s19[32],c19[32],andpr22[31],c20[32],s20[31]);


full_add fa20_32(s19[33],c19[33],andpr22[32],c20[33],s20[32]);


full_add fa20_33(s19[34],c19[34],andpr22[33],c20[34],s20[33]);


full_add fa20_34(s19[35],c19[35],andpr22[34],c20[35],s20[34]);


full_add fa20_35(s19[36],c19[36],andpr22[35],c20[36],s20[35]);


full_add fa20_36(s19[37],c19[37],andpr22[36],c20[37],s20[36]);


full_add fa20_37(s19[38],c19[38],andpr22[37],c20[38],s20[37]);


full_add fa20_38(s19[39],c19[39],andpr22[38],c20[39],s20[38]);


full_add fa20_39(s19[40],c19[40],andpr22[39],c20[40],s20[39]);


full_add fa20_40(s19[41],c19[41],andpr22[40],c20[41],s20[40]);


full_add fa20_41(s19[42],c19[42],andpr22[41],c20[42],s20[41]);


full_add fa20_42(s19[43],c19[43],andpr22[42],c20[43],s20[42]);


full_add fa20_43(s19[44],c19[44],andpr22[43],c20[44],s20[43]);


full_add fa20_44(s19[45],c19[45],andpr22[44],c20[45],s20[44]);


full_add fa20_45(s19[46],c19[46],andpr22[45],c20[46],s20[45]);


full_add fa20_46(s19[47],c19[47],andpr22[46],c20[47],s20[46]);


full_add fa20_47(s19[48],c19[48],andpr22[47],c20[48],s20[47]);


full_add fa20_48(s19[49],c19[49],andpr22[48],c20[49],s20[48]);


full_add fa20_49(s19[50],c19[50],andpr22[49],c20[50],s20[49]);


full_add fa20_50(s19[51],c19[51],andpr22[50],c20[51],s20[50]);


full_add fa20_51(s19[52],c19[52],andpr22[51],c20[52],s20[51]);


full_add fa20_52(s19[53],c19[53],andpr22[52],c20[53],s20[52]);


full_add fa20_53(s19[54],c19[54],andpr22[53],c20[54],s20[53]);


full_add fa20_54(s19[55],c19[55],andpr22[54],c20[55],s20[54]);


full_add fa20_55(s19[56],c19[56],andpr22[55],c20[56],s20[55]);


full_add fa20_56(s19[57],c19[57],andpr22[56],c20[57],s20[56]);


full_add fa20_57(s19[58],c19[58],andpr22[57],c20[58],s20[57]);


full_add fa20_58(s19[59],c19[59],andpr22[58],c20[59],s20[58]);


full_add fa20_59(s19[60],c19[60],andpr22[59],c20[60],s20[59]);


full_add fa20_60(s19[61],c19[61],andpr22[60],c20[61],s20[60]);


full_add fa20_61(s19[62],c19[62],andpr22[61],c20[62],s20[61]);


full_add fa20_62(si[20],c19[63],andpr22[62],c20[63],s20[62]);



half_adder ha21(s20[0],c20[0],c21[0],p[21]);


full_add fa21_0(s20[1],c20[1],andpr23[0],c21[1],s21[0]);


full_add fa21_1(s20[2],c20[2],andpr23[1],c21[2],s21[1]);


full_add fa21_2(s20[3],c20[3],andpr23[2],c21[3],s21[2]);


full_add fa21_3(s20[4],c20[4],andpr23[3],c21[4],s21[3]);


full_add fa21_4(s20[5],c20[5],andpr23[4],c21[5],s21[4]);


full_add fa21_5(s20[6],c20[6],andpr23[5],c21[6],s21[5]);


full_add fa21_6(s20[7],c20[7],andpr23[6],c21[7],s21[6]);


full_add fa21_7(s20[8],c20[8],andpr23[7],c21[8],s21[7]);


full_add fa21_8(s20[9],c20[9],andpr23[8],c21[9],s21[8]);


full_add fa21_9(s20[10],c20[10],andpr23[9],c21[10],s21[9]);


full_add fa21_10(s20[11],c20[11],andpr23[10],c21[11],s21[10]);


full_add fa21_11(s20[12],c20[12],andpr23[11],c21[12],s21[11]);


full_add fa21_12(s20[13],c20[13],andpr23[12],c21[13],s21[12]);


full_add fa21_13(s20[14],c20[14],andpr23[13],c21[14],s21[13]);


full_add fa21_14(s20[15],c20[15],andpr23[14],c21[15],s21[14]);


full_add fa21_15(s20[16],c20[16],andpr23[15],c21[16],s21[15]);


full_add fa21_16(s20[17],c20[17],andpr23[16],c21[17],s21[16]);


full_add fa21_17(s20[18],c20[18],andpr23[17],c21[18],s21[17]);


full_add fa21_18(s20[19],c20[19],andpr23[18],c21[19],s21[18]);


full_add fa21_19(s20[20],c20[20],andpr23[19],c21[20],s21[19]);


full_add fa21_20(s20[21],c20[21],andpr23[20],c21[21],s21[20]);


full_add fa21_21(s20[22],c20[22],andpr23[21],c21[22],s21[21]);


full_add fa21_22(s20[23],c20[23],andpr23[22],c21[23],s21[22]);


full_add fa21_23(s20[24],c20[24],andpr23[23],c21[24],s21[23]);


full_add fa21_24(s20[25],c20[25],andpr23[24],c21[25],s21[24]);


full_add fa21_25(s20[26],c20[26],andpr23[25],c21[26],s21[25]);


full_add fa21_26(s20[27],c20[27],andpr23[26],c21[27],s21[26]);


full_add fa21_27(s20[28],c20[28],andpr23[27],c21[28],s21[27]);


full_add fa21_28(s20[29],c20[29],andpr23[28],c21[29],s21[28]);


full_add fa21_29(s20[30],c20[30],andpr23[29],c21[30],s21[29]);


full_add fa21_30(s20[31],c20[31],andpr23[30],c21[31],s21[30]);


full_add fa21_31(s20[32],c20[32],andpr23[31],c21[32],s21[31]);


full_add fa21_32(s20[33],c20[33],andpr23[32],c21[33],s21[32]);


full_add fa21_33(s20[34],c20[34],andpr23[33],c21[34],s21[33]);


full_add fa21_34(s20[35],c20[35],andpr23[34],c21[35],s21[34]);


full_add fa21_35(s20[36],c20[36],andpr23[35],c21[36],s21[35]);


full_add fa21_36(s20[37],c20[37],andpr23[36],c21[37],s21[36]);


full_add fa21_37(s20[38],c20[38],andpr23[37],c21[38],s21[37]);


full_add fa21_38(s20[39],c20[39],andpr23[38],c21[39],s21[38]);


full_add fa21_39(s20[40],c20[40],andpr23[39],c21[40],s21[39]);


full_add fa21_40(s20[41],c20[41],andpr23[40],c21[41],s21[40]);


full_add fa21_41(s20[42],c20[42],andpr23[41],c21[42],s21[41]);


full_add fa21_42(s20[43],c20[43],andpr23[42],c21[43],s21[42]);


full_add fa21_43(s20[44],c20[44],andpr23[43],c21[44],s21[43]);


full_add fa21_44(s20[45],c20[45],andpr23[44],c21[45],s21[44]);


full_add fa21_45(s20[46],c20[46],andpr23[45],c21[46],s21[45]);


full_add fa21_46(s20[47],c20[47],andpr23[46],c21[47],s21[46]);


full_add fa21_47(s20[48],c20[48],andpr23[47],c21[48],s21[47]);


full_add fa21_48(s20[49],c20[49],andpr23[48],c21[49],s21[48]);


full_add fa21_49(s20[50],c20[50],andpr23[49],c21[50],s21[49]);


full_add fa21_50(s20[51],c20[51],andpr23[50],c21[51],s21[50]);


full_add fa21_51(s20[52],c20[52],andpr23[51],c21[52],s21[51]);


full_add fa21_52(s20[53],c20[53],andpr23[52],c21[53],s21[52]);


full_add fa21_53(s20[54],c20[54],andpr23[53],c21[54],s21[53]);


full_add fa21_54(s20[55],c20[55],andpr23[54],c21[55],s21[54]);


full_add fa21_55(s20[56],c20[56],andpr23[55],c21[56],s21[55]);


full_add fa21_56(s20[57],c20[57],andpr23[56],c21[57],s21[56]);


full_add fa21_57(s20[58],c20[58],andpr23[57],c21[58],s21[57]);


full_add fa21_58(s20[59],c20[59],andpr23[58],c21[59],s21[58]);


full_add fa21_59(s20[60],c20[60],andpr23[59],c21[60],s21[59]);


full_add fa21_60(s20[61],c20[61],andpr23[60],c21[61],s21[60]);


full_add fa21_61(s20[62],c20[62],andpr23[61],c21[62],s21[61]);


full_add fa21_62(si[21],c20[63],andpr23[62],c21[63],s21[62]);



half_adder ha22(s21[0],c21[0],c22[0],p[22]);


full_add fa22_0(s21[1],c21[1],andpr24[0],c22[1],s22[0]);


full_add fa22_1(s21[2],c21[2],andpr24[1],c22[2],s22[1]);


full_add fa22_2(s21[3],c21[3],andpr24[2],c22[3],s22[2]);


full_add fa22_3(s21[4],c21[4],andpr24[3],c22[4],s22[3]);


full_add fa22_4(s21[5],c21[5],andpr24[4],c22[5],s22[4]);


full_add fa22_5(s21[6],c21[6],andpr24[5],c22[6],s22[5]);


full_add fa22_6(s21[7],c21[7],andpr24[6],c22[7],s22[6]);


full_add fa22_7(s21[8],c21[8],andpr24[7],c22[8],s22[7]);


full_add fa22_8(s21[9],c21[9],andpr24[8],c22[9],s22[8]);


full_add fa22_9(s21[10],c21[10],andpr24[9],c22[10],s22[9]);


full_add fa22_10(s21[11],c21[11],andpr24[10],c22[11],s22[10]);


full_add fa22_11(s21[12],c21[12],andpr24[11],c22[12],s22[11]);


full_add fa22_12(s21[13],c21[13],andpr24[12],c22[13],s22[12]);


full_add fa22_13(s21[14],c21[14],andpr24[13],c22[14],s22[13]);


full_add fa22_14(s21[15],c21[15],andpr24[14],c22[15],s22[14]);


full_add fa22_15(s21[16],c21[16],andpr24[15],c22[16],s22[15]);


full_add fa22_16(s21[17],c21[17],andpr24[16],c22[17],s22[16]);


full_add fa22_17(s21[18],c21[18],andpr24[17],c22[18],s22[17]);


full_add fa22_18(s21[19],c21[19],andpr24[18],c22[19],s22[18]);


full_add fa22_19(s21[20],c21[20],andpr24[19],c22[20],s22[19]);


full_add fa22_20(s21[21],c21[21],andpr24[20],c22[21],s22[20]);


full_add fa22_21(s21[22],c21[22],andpr24[21],c22[22],s22[21]);


full_add fa22_22(s21[23],c21[23],andpr24[22],c22[23],s22[22]);


full_add fa22_23(s21[24],c21[24],andpr24[23],c22[24],s22[23]);


full_add fa22_24(s21[25],c21[25],andpr24[24],c22[25],s22[24]);


full_add fa22_25(s21[26],c21[26],andpr24[25],c22[26],s22[25]);


full_add fa22_26(s21[27],c21[27],andpr24[26],c22[27],s22[26]);


full_add fa22_27(s21[28],c21[28],andpr24[27],c22[28],s22[27]);


full_add fa22_28(s21[29],c21[29],andpr24[28],c22[29],s22[28]);


full_add fa22_29(s21[30],c21[30],andpr24[29],c22[30],s22[29]);


full_add fa22_30(s21[31],c21[31],andpr24[30],c22[31],s22[30]);


full_add fa22_31(s21[32],c21[32],andpr24[31],c22[32],s22[31]);


full_add fa22_32(s21[33],c21[33],andpr24[32],c22[33],s22[32]);


full_add fa22_33(s21[34],c21[34],andpr24[33],c22[34],s22[33]);


full_add fa22_34(s21[35],c21[35],andpr24[34],c22[35],s22[34]);


full_add fa22_35(s21[36],c21[36],andpr24[35],c22[36],s22[35]);


full_add fa22_36(s21[37],c21[37],andpr24[36],c22[37],s22[36]);


full_add fa22_37(s21[38],c21[38],andpr24[37],c22[38],s22[37]);


full_add fa22_38(s21[39],c21[39],andpr24[38],c22[39],s22[38]);


full_add fa22_39(s21[40],c21[40],andpr24[39],c22[40],s22[39]);


full_add fa22_40(s21[41],c21[41],andpr24[40],c22[41],s22[40]);


full_add fa22_41(s21[42],c21[42],andpr24[41],c22[42],s22[41]);


full_add fa22_42(s21[43],c21[43],andpr24[42],c22[43],s22[42]);


full_add fa22_43(s21[44],c21[44],andpr24[43],c22[44],s22[43]);


full_add fa22_44(s21[45],c21[45],andpr24[44],c22[45],s22[44]);


full_add fa22_45(s21[46],c21[46],andpr24[45],c22[46],s22[45]);


full_add fa22_46(s21[47],c21[47],andpr24[46],c22[47],s22[46]);


full_add fa22_47(s21[48],c21[48],andpr24[47],c22[48],s22[47]);


full_add fa22_48(s21[49],c21[49],andpr24[48],c22[49],s22[48]);


full_add fa22_49(s21[50],c21[50],andpr24[49],c22[50],s22[49]);


full_add fa22_50(s21[51],c21[51],andpr24[50],c22[51],s22[50]);


full_add fa22_51(s21[52],c21[52],andpr24[51],c22[52],s22[51]);


full_add fa22_52(s21[53],c21[53],andpr24[52],c22[53],s22[52]);


full_add fa22_53(s21[54],c21[54],andpr24[53],c22[54],s22[53]);


full_add fa22_54(s21[55],c21[55],andpr24[54],c22[55],s22[54]);


full_add fa22_55(s21[56],c21[56],andpr24[55],c22[56],s22[55]);


full_add fa22_56(s21[57],c21[57],andpr24[56],c22[57],s22[56]);


full_add fa22_57(s21[58],c21[58],andpr24[57],c22[58],s22[57]);


full_add fa22_58(s21[59],c21[59],andpr24[58],c22[59],s22[58]);


full_add fa22_59(s21[60],c21[60],andpr24[59],c22[60],s22[59]);


full_add fa22_60(s21[61],c21[61],andpr24[60],c22[61],s22[60]);


full_add fa22_61(s21[62],c21[62],andpr24[61],c22[62],s22[61]);


full_add fa22_62(si[22],c21[63],andpr24[62],c22[63],s22[62]);



half_adder ha23(s22[0],c22[0],c23[0],p[23]);


full_add fa23_0(s22[1],c22[1],andpr25[0],c23[1],s23[0]);


full_add fa23_1(s22[2],c22[2],andpr25[1],c23[2],s23[1]);


full_add fa23_2(s22[3],c22[3],andpr25[2],c23[3],s23[2]);


full_add fa23_3(s22[4],c22[4],andpr25[3],c23[4],s23[3]);


full_add fa23_4(s22[5],c22[5],andpr25[4],c23[5],s23[4]);


full_add fa23_5(s22[6],c22[6],andpr25[5],c23[6],s23[5]);


full_add fa23_6(s22[7],c22[7],andpr25[6],c23[7],s23[6]);


full_add fa23_7(s22[8],c22[8],andpr25[7],c23[8],s23[7]);


full_add fa23_8(s22[9],c22[9],andpr25[8],c23[9],s23[8]);


full_add fa23_9(s22[10],c22[10],andpr25[9],c23[10],s23[9]);


full_add fa23_10(s22[11],c22[11],andpr25[10],c23[11],s23[10]);


full_add fa23_11(s22[12],c22[12],andpr25[11],c23[12],s23[11]);


full_add fa23_12(s22[13],c22[13],andpr25[12],c23[13],s23[12]);


full_add fa23_13(s22[14],c22[14],andpr25[13],c23[14],s23[13]);


full_add fa23_14(s22[15],c22[15],andpr25[14],c23[15],s23[14]);


full_add fa23_15(s22[16],c22[16],andpr25[15],c23[16],s23[15]);


full_add fa23_16(s22[17],c22[17],andpr25[16],c23[17],s23[16]);


full_add fa23_17(s22[18],c22[18],andpr25[17],c23[18],s23[17]);


full_add fa23_18(s22[19],c22[19],andpr25[18],c23[19],s23[18]);


full_add fa23_19(s22[20],c22[20],andpr25[19],c23[20],s23[19]);


full_add fa23_20(s22[21],c22[21],andpr25[20],c23[21],s23[20]);


full_add fa23_21(s22[22],c22[22],andpr25[21],c23[22],s23[21]);


full_add fa23_22(s22[23],c22[23],andpr25[22],c23[23],s23[22]);


full_add fa23_23(s22[24],c22[24],andpr25[23],c23[24],s23[23]);


full_add fa23_24(s22[25],c22[25],andpr25[24],c23[25],s23[24]);


full_add fa23_25(s22[26],c22[26],andpr25[25],c23[26],s23[25]);


full_add fa23_26(s22[27],c22[27],andpr25[26],c23[27],s23[26]);


full_add fa23_27(s22[28],c22[28],andpr25[27],c23[28],s23[27]);


full_add fa23_28(s22[29],c22[29],andpr25[28],c23[29],s23[28]);


full_add fa23_29(s22[30],c22[30],andpr25[29],c23[30],s23[29]);


full_add fa23_30(s22[31],c22[31],andpr25[30],c23[31],s23[30]);


full_add fa23_31(s22[32],c22[32],andpr25[31],c23[32],s23[31]);


full_add fa23_32(s22[33],c22[33],andpr25[32],c23[33],s23[32]);


full_add fa23_33(s22[34],c22[34],andpr25[33],c23[34],s23[33]);


full_add fa23_34(s22[35],c22[35],andpr25[34],c23[35],s23[34]);


full_add fa23_35(s22[36],c22[36],andpr25[35],c23[36],s23[35]);


full_add fa23_36(s22[37],c22[37],andpr25[36],c23[37],s23[36]);


full_add fa23_37(s22[38],c22[38],andpr25[37],c23[38],s23[37]);


full_add fa23_38(s22[39],c22[39],andpr25[38],c23[39],s23[38]);


full_add fa23_39(s22[40],c22[40],andpr25[39],c23[40],s23[39]);


full_add fa23_40(s22[41],c22[41],andpr25[40],c23[41],s23[40]);


full_add fa23_41(s22[42],c22[42],andpr25[41],c23[42],s23[41]);


full_add fa23_42(s22[43],c22[43],andpr25[42],c23[43],s23[42]);


full_add fa23_43(s22[44],c22[44],andpr25[43],c23[44],s23[43]);


full_add fa23_44(s22[45],c22[45],andpr25[44],c23[45],s23[44]);


full_add fa23_45(s22[46],c22[46],andpr25[45],c23[46],s23[45]);


full_add fa23_46(s22[47],c22[47],andpr25[46],c23[47],s23[46]);


full_add fa23_47(s22[48],c22[48],andpr25[47],c23[48],s23[47]);


full_add fa23_48(s22[49],c22[49],andpr25[48],c23[49],s23[48]);


full_add fa23_49(s22[50],c22[50],andpr25[49],c23[50],s23[49]);


full_add fa23_50(s22[51],c22[51],andpr25[50],c23[51],s23[50]);


full_add fa23_51(s22[52],c22[52],andpr25[51],c23[52],s23[51]);


full_add fa23_52(s22[53],c22[53],andpr25[52],c23[53],s23[52]);


full_add fa23_53(s22[54],c22[54],andpr25[53],c23[54],s23[53]);


full_add fa23_54(s22[55],c22[55],andpr25[54],c23[55],s23[54]);


full_add fa23_55(s22[56],c22[56],andpr25[55],c23[56],s23[55]);


full_add fa23_56(s22[57],c22[57],andpr25[56],c23[57],s23[56]);


full_add fa23_57(s22[58],c22[58],andpr25[57],c23[58],s23[57]);


full_add fa23_58(s22[59],c22[59],andpr25[58],c23[59],s23[58]);


full_add fa23_59(s22[60],c22[60],andpr25[59],c23[60],s23[59]);


full_add fa23_60(s22[61],c22[61],andpr25[60],c23[61],s23[60]);


full_add fa23_61(s22[62],c22[62],andpr25[61],c23[62],s23[61]);


full_add fa23_62(si[23],c22[63],andpr25[62],c23[63],s23[62]);



half_adder ha24(s23[0],c23[0],c24[0],p[24]);


full_add fa24_0(s23[1],c23[1],andpr26[0],c24[1],s24[0]);


full_add fa24_1(s23[2],c23[2],andpr26[1],c24[2],s24[1]);


full_add fa24_2(s23[3],c23[3],andpr26[2],c24[3],s24[2]);


full_add fa24_3(s23[4],c23[4],andpr26[3],c24[4],s24[3]);


full_add fa24_4(s23[5],c23[5],andpr26[4],c24[5],s24[4]);


full_add fa24_5(s23[6],c23[6],andpr26[5],c24[6],s24[5]);


full_add fa24_6(s23[7],c23[7],andpr26[6],c24[7],s24[6]);


full_add fa24_7(s23[8],c23[8],andpr26[7],c24[8],s24[7]);


full_add fa24_8(s23[9],c23[9],andpr26[8],c24[9],s24[8]);


full_add fa24_9(s23[10],c23[10],andpr26[9],c24[10],s24[9]);


full_add fa24_10(s23[11],c23[11],andpr26[10],c24[11],s24[10]);


full_add fa24_11(s23[12],c23[12],andpr26[11],c24[12],s24[11]);


full_add fa24_12(s23[13],c23[13],andpr26[12],c24[13],s24[12]);


full_add fa24_13(s23[14],c23[14],andpr26[13],c24[14],s24[13]);


full_add fa24_14(s23[15],c23[15],andpr26[14],c24[15],s24[14]);


full_add fa24_15(s23[16],c23[16],andpr26[15],c24[16],s24[15]);


full_add fa24_16(s23[17],c23[17],andpr26[16],c24[17],s24[16]);


full_add fa24_17(s23[18],c23[18],andpr26[17],c24[18],s24[17]);


full_add fa24_18(s23[19],c23[19],andpr26[18],c24[19],s24[18]);


full_add fa24_19(s23[20],c23[20],andpr26[19],c24[20],s24[19]);


full_add fa24_20(s23[21],c23[21],andpr26[20],c24[21],s24[20]);


full_add fa24_21(s23[22],c23[22],andpr26[21],c24[22],s24[21]);


full_add fa24_22(s23[23],c23[23],andpr26[22],c24[23],s24[22]);


full_add fa24_23(s23[24],c23[24],andpr26[23],c24[24],s24[23]);


full_add fa24_24(s23[25],c23[25],andpr26[24],c24[25],s24[24]);


full_add fa24_25(s23[26],c23[26],andpr26[25],c24[26],s24[25]);


full_add fa24_26(s23[27],c23[27],andpr26[26],c24[27],s24[26]);


full_add fa24_27(s23[28],c23[28],andpr26[27],c24[28],s24[27]);


full_add fa24_28(s23[29],c23[29],andpr26[28],c24[29],s24[28]);


full_add fa24_29(s23[30],c23[30],andpr26[29],c24[30],s24[29]);


full_add fa24_30(s23[31],c23[31],andpr26[30],c24[31],s24[30]);


full_add fa24_31(s23[32],c23[32],andpr26[31],c24[32],s24[31]);


full_add fa24_32(s23[33],c23[33],andpr26[32],c24[33],s24[32]);


full_add fa24_33(s23[34],c23[34],andpr26[33],c24[34],s24[33]);


full_add fa24_34(s23[35],c23[35],andpr26[34],c24[35],s24[34]);


full_add fa24_35(s23[36],c23[36],andpr26[35],c24[36],s24[35]);


full_add fa24_36(s23[37],c23[37],andpr26[36],c24[37],s24[36]);


full_add fa24_37(s23[38],c23[38],andpr26[37],c24[38],s24[37]);


full_add fa24_38(s23[39],c23[39],andpr26[38],c24[39],s24[38]);


full_add fa24_39(s23[40],c23[40],andpr26[39],c24[40],s24[39]);


full_add fa24_40(s23[41],c23[41],andpr26[40],c24[41],s24[40]);


full_add fa24_41(s23[42],c23[42],andpr26[41],c24[42],s24[41]);


full_add fa24_42(s23[43],c23[43],andpr26[42],c24[43],s24[42]);


full_add fa24_43(s23[44],c23[44],andpr26[43],c24[44],s24[43]);


full_add fa24_44(s23[45],c23[45],andpr26[44],c24[45],s24[44]);


full_add fa24_45(s23[46],c23[46],andpr26[45],c24[46],s24[45]);


full_add fa24_46(s23[47],c23[47],andpr26[46],c24[47],s24[46]);


full_add fa24_47(s23[48],c23[48],andpr26[47],c24[48],s24[47]);


full_add fa24_48(s23[49],c23[49],andpr26[48],c24[49],s24[48]);


full_add fa24_49(s23[50],c23[50],andpr26[49],c24[50],s24[49]);


full_add fa24_50(s23[51],c23[51],andpr26[50],c24[51],s24[50]);


full_add fa24_51(s23[52],c23[52],andpr26[51],c24[52],s24[51]);


full_add fa24_52(s23[53],c23[53],andpr26[52],c24[53],s24[52]);


full_add fa24_53(s23[54],c23[54],andpr26[53],c24[54],s24[53]);


full_add fa24_54(s23[55],c23[55],andpr26[54],c24[55],s24[54]);


full_add fa24_55(s23[56],c23[56],andpr26[55],c24[56],s24[55]);


full_add fa24_56(s23[57],c23[57],andpr26[56],c24[57],s24[56]);


full_add fa24_57(s23[58],c23[58],andpr26[57],c24[58],s24[57]);


full_add fa24_58(s23[59],c23[59],andpr26[58],c24[59],s24[58]);


full_add fa24_59(s23[60],c23[60],andpr26[59],c24[60],s24[59]);


full_add fa24_60(s23[61],c23[61],andpr26[60],c24[61],s24[60]);


full_add fa24_61(s23[62],c23[62],andpr26[61],c24[62],s24[61]);


full_add fa24_62(si[24],c23[63],andpr26[62],c24[63],s24[62]);



half_adder ha25(s24[0],c24[0],c25[0],p[25]);


full_add fa25_0(s24[1],c24[1],andpr27[0],c25[1],s25[0]);


full_add fa25_1(s24[2],c24[2],andpr27[1],c25[2],s25[1]);


full_add fa25_2(s24[3],c24[3],andpr27[2],c25[3],s25[2]);


full_add fa25_3(s24[4],c24[4],andpr27[3],c25[4],s25[3]);


full_add fa25_4(s24[5],c24[5],andpr27[4],c25[5],s25[4]);


full_add fa25_5(s24[6],c24[6],andpr27[5],c25[6],s25[5]);


full_add fa25_6(s24[7],c24[7],andpr27[6],c25[7],s25[6]);


full_add fa25_7(s24[8],c24[8],andpr27[7],c25[8],s25[7]);


full_add fa25_8(s24[9],c24[9],andpr27[8],c25[9],s25[8]);


full_add fa25_9(s24[10],c24[10],andpr27[9],c25[10],s25[9]);


full_add fa25_10(s24[11],c24[11],andpr27[10],c25[11],s25[10]);


full_add fa25_11(s24[12],c24[12],andpr27[11],c25[12],s25[11]);


full_add fa25_12(s24[13],c24[13],andpr27[12],c25[13],s25[12]);


full_add fa25_13(s24[14],c24[14],andpr27[13],c25[14],s25[13]);


full_add fa25_14(s24[15],c24[15],andpr27[14],c25[15],s25[14]);


full_add fa25_15(s24[16],c24[16],andpr27[15],c25[16],s25[15]);


full_add fa25_16(s24[17],c24[17],andpr27[16],c25[17],s25[16]);


full_add fa25_17(s24[18],c24[18],andpr27[17],c25[18],s25[17]);


full_add fa25_18(s24[19],c24[19],andpr27[18],c25[19],s25[18]);


full_add fa25_19(s24[20],c24[20],andpr27[19],c25[20],s25[19]);


full_add fa25_20(s24[21],c24[21],andpr27[20],c25[21],s25[20]);


full_add fa25_21(s24[22],c24[22],andpr27[21],c25[22],s25[21]);


full_add fa25_22(s24[23],c24[23],andpr27[22],c25[23],s25[22]);


full_add fa25_23(s24[24],c24[24],andpr27[23],c25[24],s25[23]);


full_add fa25_24(s24[25],c24[25],andpr27[24],c25[25],s25[24]);


full_add fa25_25(s24[26],c24[26],andpr27[25],c25[26],s25[25]);


full_add fa25_26(s24[27],c24[27],andpr27[26],c25[27],s25[26]);


full_add fa25_27(s24[28],c24[28],andpr27[27],c25[28],s25[27]);


full_add fa25_28(s24[29],c24[29],andpr27[28],c25[29],s25[28]);


full_add fa25_29(s24[30],c24[30],andpr27[29],c25[30],s25[29]);


full_add fa25_30(s24[31],c24[31],andpr27[30],c25[31],s25[30]);


full_add fa25_31(s24[32],c24[32],andpr27[31],c25[32],s25[31]);


full_add fa25_32(s24[33],c24[33],andpr27[32],c25[33],s25[32]);


full_add fa25_33(s24[34],c24[34],andpr27[33],c25[34],s25[33]);


full_add fa25_34(s24[35],c24[35],andpr27[34],c25[35],s25[34]);


full_add fa25_35(s24[36],c24[36],andpr27[35],c25[36],s25[35]);


full_add fa25_36(s24[37],c24[37],andpr27[36],c25[37],s25[36]);


full_add fa25_37(s24[38],c24[38],andpr27[37],c25[38],s25[37]);


full_add fa25_38(s24[39],c24[39],andpr27[38],c25[39],s25[38]);


full_add fa25_39(s24[40],c24[40],andpr27[39],c25[40],s25[39]);


full_add fa25_40(s24[41],c24[41],andpr27[40],c25[41],s25[40]);


full_add fa25_41(s24[42],c24[42],andpr27[41],c25[42],s25[41]);


full_add fa25_42(s24[43],c24[43],andpr27[42],c25[43],s25[42]);


full_add fa25_43(s24[44],c24[44],andpr27[43],c25[44],s25[43]);


full_add fa25_44(s24[45],c24[45],andpr27[44],c25[45],s25[44]);


full_add fa25_45(s24[46],c24[46],andpr27[45],c25[46],s25[45]);


full_add fa25_46(s24[47],c24[47],andpr27[46],c25[47],s25[46]);


full_add fa25_47(s24[48],c24[48],andpr27[47],c25[48],s25[47]);


full_add fa25_48(s24[49],c24[49],andpr27[48],c25[49],s25[48]);


full_add fa25_49(s24[50],c24[50],andpr27[49],c25[50],s25[49]);


full_add fa25_50(s24[51],c24[51],andpr27[50],c25[51],s25[50]);


full_add fa25_51(s24[52],c24[52],andpr27[51],c25[52],s25[51]);


full_add fa25_52(s24[53],c24[53],andpr27[52],c25[53],s25[52]);


full_add fa25_53(s24[54],c24[54],andpr27[53],c25[54],s25[53]);


full_add fa25_54(s24[55],c24[55],andpr27[54],c25[55],s25[54]);


full_add fa25_55(s24[56],c24[56],andpr27[55],c25[56],s25[55]);


full_add fa25_56(s24[57],c24[57],andpr27[56],c25[57],s25[56]);


full_add fa25_57(s24[58],c24[58],andpr27[57],c25[58],s25[57]);


full_add fa25_58(s24[59],c24[59],andpr27[58],c25[59],s25[58]);


full_add fa25_59(s24[60],c24[60],andpr27[59],c25[60],s25[59]);


full_add fa25_60(s24[61],c24[61],andpr27[60],c25[61],s25[60]);


full_add fa25_61(s24[62],c24[62],andpr27[61],c25[62],s25[61]);


full_add fa25_62(si[25],c24[63],andpr27[62],c25[63],s25[62]);



half_adder ha26(s25[0],c25[0],c26[0],p[26]);


full_add fa26_0(s25[1],c25[1],andpr28[0],c26[1],s26[0]);


full_add fa26_1(s25[2],c25[2],andpr28[1],c26[2],s26[1]);


full_add fa26_2(s25[3],c25[3],andpr28[2],c26[3],s26[2]);


full_add fa26_3(s25[4],c25[4],andpr28[3],c26[4],s26[3]);


full_add fa26_4(s25[5],c25[5],andpr28[4],c26[5],s26[4]);


full_add fa26_5(s25[6],c25[6],andpr28[5],c26[6],s26[5]);


full_add fa26_6(s25[7],c25[7],andpr28[6],c26[7],s26[6]);


full_add fa26_7(s25[8],c25[8],andpr28[7],c26[8],s26[7]);


full_add fa26_8(s25[9],c25[9],andpr28[8],c26[9],s26[8]);


full_add fa26_9(s25[10],c25[10],andpr28[9],c26[10],s26[9]);


full_add fa26_10(s25[11],c25[11],andpr28[10],c26[11],s26[10]);


full_add fa26_11(s25[12],c25[12],andpr28[11],c26[12],s26[11]);


full_add fa26_12(s25[13],c25[13],andpr28[12],c26[13],s26[12]);


full_add fa26_13(s25[14],c25[14],andpr28[13],c26[14],s26[13]);


full_add fa26_14(s25[15],c25[15],andpr28[14],c26[15],s26[14]);


full_add fa26_15(s25[16],c25[16],andpr28[15],c26[16],s26[15]);


full_add fa26_16(s25[17],c25[17],andpr28[16],c26[17],s26[16]);


full_add fa26_17(s25[18],c25[18],andpr28[17],c26[18],s26[17]);


full_add fa26_18(s25[19],c25[19],andpr28[18],c26[19],s26[18]);


full_add fa26_19(s25[20],c25[20],andpr28[19],c26[20],s26[19]);


full_add fa26_20(s25[21],c25[21],andpr28[20],c26[21],s26[20]);


full_add fa26_21(s25[22],c25[22],andpr28[21],c26[22],s26[21]);


full_add fa26_22(s25[23],c25[23],andpr28[22],c26[23],s26[22]);


full_add fa26_23(s25[24],c25[24],andpr28[23],c26[24],s26[23]);


full_add fa26_24(s25[25],c25[25],andpr28[24],c26[25],s26[24]);


full_add fa26_25(s25[26],c25[26],andpr28[25],c26[26],s26[25]);


full_add fa26_26(s25[27],c25[27],andpr28[26],c26[27],s26[26]);


full_add fa26_27(s25[28],c25[28],andpr28[27],c26[28],s26[27]);


full_add fa26_28(s25[29],c25[29],andpr28[28],c26[29],s26[28]);


full_add fa26_29(s25[30],c25[30],andpr28[29],c26[30],s26[29]);


full_add fa26_30(s25[31],c25[31],andpr28[30],c26[31],s26[30]);


full_add fa26_31(s25[32],c25[32],andpr28[31],c26[32],s26[31]);


full_add fa26_32(s25[33],c25[33],andpr28[32],c26[33],s26[32]);


full_add fa26_33(s25[34],c25[34],andpr28[33],c26[34],s26[33]);


full_add fa26_34(s25[35],c25[35],andpr28[34],c26[35],s26[34]);


full_add fa26_35(s25[36],c25[36],andpr28[35],c26[36],s26[35]);


full_add fa26_36(s25[37],c25[37],andpr28[36],c26[37],s26[36]);


full_add fa26_37(s25[38],c25[38],andpr28[37],c26[38],s26[37]);


full_add fa26_38(s25[39],c25[39],andpr28[38],c26[39],s26[38]);


full_add fa26_39(s25[40],c25[40],andpr28[39],c26[40],s26[39]);


full_add fa26_40(s25[41],c25[41],andpr28[40],c26[41],s26[40]);


full_add fa26_41(s25[42],c25[42],andpr28[41],c26[42],s26[41]);


full_add fa26_42(s25[43],c25[43],andpr28[42],c26[43],s26[42]);


full_add fa26_43(s25[44],c25[44],andpr28[43],c26[44],s26[43]);


full_add fa26_44(s25[45],c25[45],andpr28[44],c26[45],s26[44]);


full_add fa26_45(s25[46],c25[46],andpr28[45],c26[46],s26[45]);


full_add fa26_46(s25[47],c25[47],andpr28[46],c26[47],s26[46]);


full_add fa26_47(s25[48],c25[48],andpr28[47],c26[48],s26[47]);


full_add fa26_48(s25[49],c25[49],andpr28[48],c26[49],s26[48]);


full_add fa26_49(s25[50],c25[50],andpr28[49],c26[50],s26[49]);


full_add fa26_50(s25[51],c25[51],andpr28[50],c26[51],s26[50]);


full_add fa26_51(s25[52],c25[52],andpr28[51],c26[52],s26[51]);


full_add fa26_52(s25[53],c25[53],andpr28[52],c26[53],s26[52]);


full_add fa26_53(s25[54],c25[54],andpr28[53],c26[54],s26[53]);


full_add fa26_54(s25[55],c25[55],andpr28[54],c26[55],s26[54]);


full_add fa26_55(s25[56],c25[56],andpr28[55],c26[56],s26[55]);


full_add fa26_56(s25[57],c25[57],andpr28[56],c26[57],s26[56]);


full_add fa26_57(s25[58],c25[58],andpr28[57],c26[58],s26[57]);


full_add fa26_58(s25[59],c25[59],andpr28[58],c26[59],s26[58]);


full_add fa26_59(s25[60],c25[60],andpr28[59],c26[60],s26[59]);


full_add fa26_60(s25[61],c25[61],andpr28[60],c26[61],s26[60]);


full_add fa26_61(s25[62],c25[62],andpr28[61],c26[62],s26[61]);


full_add fa26_62(si[26],c25[63],andpr28[62],c26[63],s26[62]);



half_adder ha27(s26[0],c26[0],c27[0],p[27]);


full_add fa27_0(s26[1],c26[1],andpr29[0],c27[1],s27[0]);


full_add fa27_1(s26[2],c26[2],andpr29[1],c27[2],s27[1]);


full_add fa27_2(s26[3],c26[3],andpr29[2],c27[3],s27[2]);


full_add fa27_3(s26[4],c26[4],andpr29[3],c27[4],s27[3]);


full_add fa27_4(s26[5],c26[5],andpr29[4],c27[5],s27[4]);


full_add fa27_5(s26[6],c26[6],andpr29[5],c27[6],s27[5]);


full_add fa27_6(s26[7],c26[7],andpr29[6],c27[7],s27[6]);


full_add fa27_7(s26[8],c26[8],andpr29[7],c27[8],s27[7]);


full_add fa27_8(s26[9],c26[9],andpr29[8],c27[9],s27[8]);


full_add fa27_9(s26[10],c26[10],andpr29[9],c27[10],s27[9]);


full_add fa27_10(s26[11],c26[11],andpr29[10],c27[11],s27[10]);


full_add fa27_11(s26[12],c26[12],andpr29[11],c27[12],s27[11]);


full_add fa27_12(s26[13],c26[13],andpr29[12],c27[13],s27[12]);


full_add fa27_13(s26[14],c26[14],andpr29[13],c27[14],s27[13]);


full_add fa27_14(s26[15],c26[15],andpr29[14],c27[15],s27[14]);


full_add fa27_15(s26[16],c26[16],andpr29[15],c27[16],s27[15]);


full_add fa27_16(s26[17],c26[17],andpr29[16],c27[17],s27[16]);


full_add fa27_17(s26[18],c26[18],andpr29[17],c27[18],s27[17]);


full_add fa27_18(s26[19],c26[19],andpr29[18],c27[19],s27[18]);


full_add fa27_19(s26[20],c26[20],andpr29[19],c27[20],s27[19]);


full_add fa27_20(s26[21],c26[21],andpr29[20],c27[21],s27[20]);


full_add fa27_21(s26[22],c26[22],andpr29[21],c27[22],s27[21]);


full_add fa27_22(s26[23],c26[23],andpr29[22],c27[23],s27[22]);


full_add fa27_23(s26[24],c26[24],andpr29[23],c27[24],s27[23]);


full_add fa27_24(s26[25],c26[25],andpr29[24],c27[25],s27[24]);


full_add fa27_25(s26[26],c26[26],andpr29[25],c27[26],s27[25]);


full_add fa27_26(s26[27],c26[27],andpr29[26],c27[27],s27[26]);


full_add fa27_27(s26[28],c26[28],andpr29[27],c27[28],s27[27]);


full_add fa27_28(s26[29],c26[29],andpr29[28],c27[29],s27[28]);


full_add fa27_29(s26[30],c26[30],andpr29[29],c27[30],s27[29]);


full_add fa27_30(s26[31],c26[31],andpr29[30],c27[31],s27[30]);


full_add fa27_31(s26[32],c26[32],andpr29[31],c27[32],s27[31]);


full_add fa27_32(s26[33],c26[33],andpr29[32],c27[33],s27[32]);


full_add fa27_33(s26[34],c26[34],andpr29[33],c27[34],s27[33]);


full_add fa27_34(s26[35],c26[35],andpr29[34],c27[35],s27[34]);


full_add fa27_35(s26[36],c26[36],andpr29[35],c27[36],s27[35]);


full_add fa27_36(s26[37],c26[37],andpr29[36],c27[37],s27[36]);


full_add fa27_37(s26[38],c26[38],andpr29[37],c27[38],s27[37]);


full_add fa27_38(s26[39],c26[39],andpr29[38],c27[39],s27[38]);


full_add fa27_39(s26[40],c26[40],andpr29[39],c27[40],s27[39]);


full_add fa27_40(s26[41],c26[41],andpr29[40],c27[41],s27[40]);


full_add fa27_41(s26[42],c26[42],andpr29[41],c27[42],s27[41]);


full_add fa27_42(s26[43],c26[43],andpr29[42],c27[43],s27[42]);


full_add fa27_43(s26[44],c26[44],andpr29[43],c27[44],s27[43]);


full_add fa27_44(s26[45],c26[45],andpr29[44],c27[45],s27[44]);


full_add fa27_45(s26[46],c26[46],andpr29[45],c27[46],s27[45]);


full_add fa27_46(s26[47],c26[47],andpr29[46],c27[47],s27[46]);


full_add fa27_47(s26[48],c26[48],andpr29[47],c27[48],s27[47]);


full_add fa27_48(s26[49],c26[49],andpr29[48],c27[49],s27[48]);


full_add fa27_49(s26[50],c26[50],andpr29[49],c27[50],s27[49]);


full_add fa27_50(s26[51],c26[51],andpr29[50],c27[51],s27[50]);


full_add fa27_51(s26[52],c26[52],andpr29[51],c27[52],s27[51]);


full_add fa27_52(s26[53],c26[53],andpr29[52],c27[53],s27[52]);


full_add fa27_53(s26[54],c26[54],andpr29[53],c27[54],s27[53]);


full_add fa27_54(s26[55],c26[55],andpr29[54],c27[55],s27[54]);


full_add fa27_55(s26[56],c26[56],andpr29[55],c27[56],s27[55]);


full_add fa27_56(s26[57],c26[57],andpr29[56],c27[57],s27[56]);


full_add fa27_57(s26[58],c26[58],andpr29[57],c27[58],s27[57]);


full_add fa27_58(s26[59],c26[59],andpr29[58],c27[59],s27[58]);


full_add fa27_59(s26[60],c26[60],andpr29[59],c27[60],s27[59]);


full_add fa27_60(s26[61],c26[61],andpr29[60],c27[61],s27[60]);


full_add fa27_61(s26[62],c26[62],andpr29[61],c27[62],s27[61]);


full_add fa27_62(si[27],c26[63],andpr29[62],c27[63],s27[62]);



half_adder ha28(s27[0],c27[0],c28[0],p[28]);


full_add fa28_0(s27[1],c27[1],andpr30[0],c28[1],s28[0]);


full_add fa28_1(s27[2],c27[2],andpr30[1],c28[2],s28[1]);


full_add fa28_2(s27[3],c27[3],andpr30[2],c28[3],s28[2]);


full_add fa28_3(s27[4],c27[4],andpr30[3],c28[4],s28[3]);


full_add fa28_4(s27[5],c27[5],andpr30[4],c28[5],s28[4]);


full_add fa28_5(s27[6],c27[6],andpr30[5],c28[6],s28[5]);


full_add fa28_6(s27[7],c27[7],andpr30[6],c28[7],s28[6]);


full_add fa28_7(s27[8],c27[8],andpr30[7],c28[8],s28[7]);


full_add fa28_8(s27[9],c27[9],andpr30[8],c28[9],s28[8]);


full_add fa28_9(s27[10],c27[10],andpr30[9],c28[10],s28[9]);


full_add fa28_10(s27[11],c27[11],andpr30[10],c28[11],s28[10]);


full_add fa28_11(s27[12],c27[12],andpr30[11],c28[12],s28[11]);


full_add fa28_12(s27[13],c27[13],andpr30[12],c28[13],s28[12]);


full_add fa28_13(s27[14],c27[14],andpr30[13],c28[14],s28[13]);


full_add fa28_14(s27[15],c27[15],andpr30[14],c28[15],s28[14]);


full_add fa28_15(s27[16],c27[16],andpr30[15],c28[16],s28[15]);


full_add fa28_16(s27[17],c27[17],andpr30[16],c28[17],s28[16]);


full_add fa28_17(s27[18],c27[18],andpr30[17],c28[18],s28[17]);


full_add fa28_18(s27[19],c27[19],andpr30[18],c28[19],s28[18]);


full_add fa28_19(s27[20],c27[20],andpr30[19],c28[20],s28[19]);


full_add fa28_20(s27[21],c27[21],andpr30[20],c28[21],s28[20]);


full_add fa28_21(s27[22],c27[22],andpr30[21],c28[22],s28[21]);


full_add fa28_22(s27[23],c27[23],andpr30[22],c28[23],s28[22]);


full_add fa28_23(s27[24],c27[24],andpr30[23],c28[24],s28[23]);


full_add fa28_24(s27[25],c27[25],andpr30[24],c28[25],s28[24]);


full_add fa28_25(s27[26],c27[26],andpr30[25],c28[26],s28[25]);


full_add fa28_26(s27[27],c27[27],andpr30[26],c28[27],s28[26]);


full_add fa28_27(s27[28],c27[28],andpr30[27],c28[28],s28[27]);


full_add fa28_28(s27[29],c27[29],andpr30[28],c28[29],s28[28]);


full_add fa28_29(s27[30],c27[30],andpr30[29],c28[30],s28[29]);


full_add fa28_30(s27[31],c27[31],andpr30[30],c28[31],s28[30]);


full_add fa28_31(s27[32],c27[32],andpr30[31],c28[32],s28[31]);


full_add fa28_32(s27[33],c27[33],andpr30[32],c28[33],s28[32]);


full_add fa28_33(s27[34],c27[34],andpr30[33],c28[34],s28[33]);


full_add fa28_34(s27[35],c27[35],andpr30[34],c28[35],s28[34]);


full_add fa28_35(s27[36],c27[36],andpr30[35],c28[36],s28[35]);


full_add fa28_36(s27[37],c27[37],andpr30[36],c28[37],s28[36]);


full_add fa28_37(s27[38],c27[38],andpr30[37],c28[38],s28[37]);


full_add fa28_38(s27[39],c27[39],andpr30[38],c28[39],s28[38]);


full_add fa28_39(s27[40],c27[40],andpr30[39],c28[40],s28[39]);


full_add fa28_40(s27[41],c27[41],andpr30[40],c28[41],s28[40]);


full_add fa28_41(s27[42],c27[42],andpr30[41],c28[42],s28[41]);


full_add fa28_42(s27[43],c27[43],andpr30[42],c28[43],s28[42]);


full_add fa28_43(s27[44],c27[44],andpr30[43],c28[44],s28[43]);


full_add fa28_44(s27[45],c27[45],andpr30[44],c28[45],s28[44]);


full_add fa28_45(s27[46],c27[46],andpr30[45],c28[46],s28[45]);


full_add fa28_46(s27[47],c27[47],andpr30[46],c28[47],s28[46]);


full_add fa28_47(s27[48],c27[48],andpr30[47],c28[48],s28[47]);


full_add fa28_48(s27[49],c27[49],andpr30[48],c28[49],s28[48]);


full_add fa28_49(s27[50],c27[50],andpr30[49],c28[50],s28[49]);


full_add fa28_50(s27[51],c27[51],andpr30[50],c28[51],s28[50]);


full_add fa28_51(s27[52],c27[52],andpr30[51],c28[52],s28[51]);


full_add fa28_52(s27[53],c27[53],andpr30[52],c28[53],s28[52]);


full_add fa28_53(s27[54],c27[54],andpr30[53],c28[54],s28[53]);


full_add fa28_54(s27[55],c27[55],andpr30[54],c28[55],s28[54]);


full_add fa28_55(s27[56],c27[56],andpr30[55],c28[56],s28[55]);


full_add fa28_56(s27[57],c27[57],andpr30[56],c28[57],s28[56]);


full_add fa28_57(s27[58],c27[58],andpr30[57],c28[58],s28[57]);


full_add fa28_58(s27[59],c27[59],andpr30[58],c28[59],s28[58]);


full_add fa28_59(s27[60],c27[60],andpr30[59],c28[60],s28[59]);


full_add fa28_60(s27[61],c27[61],andpr30[60],c28[61],s28[60]);


full_add fa28_61(s27[62],c27[62],andpr30[61],c28[62],s28[61]);


full_add fa28_62(si[28],c27[63],andpr30[62],c28[63],s28[62]);



half_adder ha29(s28[0],c28[0],c29[0],p[29]);


full_add fa29_0(s28[1],c28[1],andpr31[0],c29[1],s29[0]);


full_add fa29_1(s28[2],c28[2],andpr31[1],c29[2],s29[1]);


full_add fa29_2(s28[3],c28[3],andpr31[2],c29[3],s29[2]);


full_add fa29_3(s28[4],c28[4],andpr31[3],c29[4],s29[3]);


full_add fa29_4(s28[5],c28[5],andpr31[4],c29[5],s29[4]);


full_add fa29_5(s28[6],c28[6],andpr31[5],c29[6],s29[5]);


full_add fa29_6(s28[7],c28[7],andpr31[6],c29[7],s29[6]);


full_add fa29_7(s28[8],c28[8],andpr31[7],c29[8],s29[7]);


full_add fa29_8(s28[9],c28[9],andpr31[8],c29[9],s29[8]);


full_add fa29_9(s28[10],c28[10],andpr31[9],c29[10],s29[9]);


full_add fa29_10(s28[11],c28[11],andpr31[10],c29[11],s29[10]);


full_add fa29_11(s28[12],c28[12],andpr31[11],c29[12],s29[11]);


full_add fa29_12(s28[13],c28[13],andpr31[12],c29[13],s29[12]);


full_add fa29_13(s28[14],c28[14],andpr31[13],c29[14],s29[13]);


full_add fa29_14(s28[15],c28[15],andpr31[14],c29[15],s29[14]);


full_add fa29_15(s28[16],c28[16],andpr31[15],c29[16],s29[15]);


full_add fa29_16(s28[17],c28[17],andpr31[16],c29[17],s29[16]);


full_add fa29_17(s28[18],c28[18],andpr31[17],c29[18],s29[17]);


full_add fa29_18(s28[19],c28[19],andpr31[18],c29[19],s29[18]);


full_add fa29_19(s28[20],c28[20],andpr31[19],c29[20],s29[19]);


full_add fa29_20(s28[21],c28[21],andpr31[20],c29[21],s29[20]);


full_add fa29_21(s28[22],c28[22],andpr31[21],c29[22],s29[21]);


full_add fa29_22(s28[23],c28[23],andpr31[22],c29[23],s29[22]);


full_add fa29_23(s28[24],c28[24],andpr31[23],c29[24],s29[23]);


full_add fa29_24(s28[25],c28[25],andpr31[24],c29[25],s29[24]);


full_add fa29_25(s28[26],c28[26],andpr31[25],c29[26],s29[25]);


full_add fa29_26(s28[27],c28[27],andpr31[26],c29[27],s29[26]);


full_add fa29_27(s28[28],c28[28],andpr31[27],c29[28],s29[27]);


full_add fa29_28(s28[29],c28[29],andpr31[28],c29[29],s29[28]);


full_add fa29_29(s28[30],c28[30],andpr31[29],c29[30],s29[29]);


full_add fa29_30(s28[31],c28[31],andpr31[30],c29[31],s29[30]);


full_add fa29_31(s28[32],c28[32],andpr31[31],c29[32],s29[31]);


full_add fa29_32(s28[33],c28[33],andpr31[32],c29[33],s29[32]);


full_add fa29_33(s28[34],c28[34],andpr31[33],c29[34],s29[33]);


full_add fa29_34(s28[35],c28[35],andpr31[34],c29[35],s29[34]);


full_add fa29_35(s28[36],c28[36],andpr31[35],c29[36],s29[35]);


full_add fa29_36(s28[37],c28[37],andpr31[36],c29[37],s29[36]);


full_add fa29_37(s28[38],c28[38],andpr31[37],c29[38],s29[37]);


full_add fa29_38(s28[39],c28[39],andpr31[38],c29[39],s29[38]);


full_add fa29_39(s28[40],c28[40],andpr31[39],c29[40],s29[39]);


full_add fa29_40(s28[41],c28[41],andpr31[40],c29[41],s29[40]);


full_add fa29_41(s28[42],c28[42],andpr31[41],c29[42],s29[41]);


full_add fa29_42(s28[43],c28[43],andpr31[42],c29[43],s29[42]);


full_add fa29_43(s28[44],c28[44],andpr31[43],c29[44],s29[43]);


full_add fa29_44(s28[45],c28[45],andpr31[44],c29[45],s29[44]);


full_add fa29_45(s28[46],c28[46],andpr31[45],c29[46],s29[45]);


full_add fa29_46(s28[47],c28[47],andpr31[46],c29[47],s29[46]);


full_add fa29_47(s28[48],c28[48],andpr31[47],c29[48],s29[47]);


full_add fa29_48(s28[49],c28[49],andpr31[48],c29[49],s29[48]);


full_add fa29_49(s28[50],c28[50],andpr31[49],c29[50],s29[49]);


full_add fa29_50(s28[51],c28[51],andpr31[50],c29[51],s29[50]);


full_add fa29_51(s28[52],c28[52],andpr31[51],c29[52],s29[51]);


full_add fa29_52(s28[53],c28[53],andpr31[52],c29[53],s29[52]);


full_add fa29_53(s28[54],c28[54],andpr31[53],c29[54],s29[53]);


full_add fa29_54(s28[55],c28[55],andpr31[54],c29[55],s29[54]);


full_add fa29_55(s28[56],c28[56],andpr31[55],c29[56],s29[55]);


full_add fa29_56(s28[57],c28[57],andpr31[56],c29[57],s29[56]);


full_add fa29_57(s28[58],c28[58],andpr31[57],c29[58],s29[57]);


full_add fa29_58(s28[59],c28[59],andpr31[58],c29[59],s29[58]);


full_add fa29_59(s28[60],c28[60],andpr31[59],c29[60],s29[59]);


full_add fa29_60(s28[61],c28[61],andpr31[60],c29[61],s29[60]);


full_add fa29_61(s28[62],c28[62],andpr31[61],c29[62],s29[61]);


full_add fa29_62(si[29],c28[63],andpr31[62],c29[63],s29[62]);



half_adder ha30(s29[0],c29[0],c30[0],p[30]);


full_add fa30_0(s29[1],c29[1],andpr32[0],c30[1],s30[0]);


full_add fa30_1(s29[2],c29[2],andpr32[1],c30[2],s30[1]);


full_add fa30_2(s29[3],c29[3],andpr32[2],c30[3],s30[2]);


full_add fa30_3(s29[4],c29[4],andpr32[3],c30[4],s30[3]);


full_add fa30_4(s29[5],c29[5],andpr32[4],c30[5],s30[4]);


full_add fa30_5(s29[6],c29[6],andpr32[5],c30[6],s30[5]);


full_add fa30_6(s29[7],c29[7],andpr32[6],c30[7],s30[6]);


full_add fa30_7(s29[8],c29[8],andpr32[7],c30[8],s30[7]);


full_add fa30_8(s29[9],c29[9],andpr32[8],c30[9],s30[8]);


full_add fa30_9(s29[10],c29[10],andpr32[9],c30[10],s30[9]);


full_add fa30_10(s29[11],c29[11],andpr32[10],c30[11],s30[10]);


full_add fa30_11(s29[12],c29[12],andpr32[11],c30[12],s30[11]);


full_add fa30_12(s29[13],c29[13],andpr32[12],c30[13],s30[12]);


full_add fa30_13(s29[14],c29[14],andpr32[13],c30[14],s30[13]);


full_add fa30_14(s29[15],c29[15],andpr32[14],c30[15],s30[14]);


full_add fa30_15(s29[16],c29[16],andpr32[15],c30[16],s30[15]);


full_add fa30_16(s29[17],c29[17],andpr32[16],c30[17],s30[16]);


full_add fa30_17(s29[18],c29[18],andpr32[17],c30[18],s30[17]);


full_add fa30_18(s29[19],c29[19],andpr32[18],c30[19],s30[18]);


full_add fa30_19(s29[20],c29[20],andpr32[19],c30[20],s30[19]);


full_add fa30_20(s29[21],c29[21],andpr32[20],c30[21],s30[20]);


full_add fa30_21(s29[22],c29[22],andpr32[21],c30[22],s30[21]);


full_add fa30_22(s29[23],c29[23],andpr32[22],c30[23],s30[22]);


full_add fa30_23(s29[24],c29[24],andpr32[23],c30[24],s30[23]);


full_add fa30_24(s29[25],c29[25],andpr32[24],c30[25],s30[24]);


full_add fa30_25(s29[26],c29[26],andpr32[25],c30[26],s30[25]);


full_add fa30_26(s29[27],c29[27],andpr32[26],c30[27],s30[26]);


full_add fa30_27(s29[28],c29[28],andpr32[27],c30[28],s30[27]);


full_add fa30_28(s29[29],c29[29],andpr32[28],c30[29],s30[28]);


full_add fa30_29(s29[30],c29[30],andpr32[29],c30[30],s30[29]);


full_add fa30_30(s29[31],c29[31],andpr32[30],c30[31],s30[30]);


full_add fa30_31(s29[32],c29[32],andpr32[31],c30[32],s30[31]);


full_add fa30_32(s29[33],c29[33],andpr32[32],c30[33],s30[32]);


full_add fa30_33(s29[34],c29[34],andpr32[33],c30[34],s30[33]);


full_add fa30_34(s29[35],c29[35],andpr32[34],c30[35],s30[34]);


full_add fa30_35(s29[36],c29[36],andpr32[35],c30[36],s30[35]);


full_add fa30_36(s29[37],c29[37],andpr32[36],c30[37],s30[36]);


full_add fa30_37(s29[38],c29[38],andpr32[37],c30[38],s30[37]);


full_add fa30_38(s29[39],c29[39],andpr32[38],c30[39],s30[38]);


full_add fa30_39(s29[40],c29[40],andpr32[39],c30[40],s30[39]);


full_add fa30_40(s29[41],c29[41],andpr32[40],c30[41],s30[40]);


full_add fa30_41(s29[42],c29[42],andpr32[41],c30[42],s30[41]);


full_add fa30_42(s29[43],c29[43],andpr32[42],c30[43],s30[42]);


full_add fa30_43(s29[44],c29[44],andpr32[43],c30[44],s30[43]);


full_add fa30_44(s29[45],c29[45],andpr32[44],c30[45],s30[44]);


full_add fa30_45(s29[46],c29[46],andpr32[45],c30[46],s30[45]);


full_add fa30_46(s29[47],c29[47],andpr32[46],c30[47],s30[46]);


full_add fa30_47(s29[48],c29[48],andpr32[47],c30[48],s30[47]);


full_add fa30_48(s29[49],c29[49],andpr32[48],c30[49],s30[48]);


full_add fa30_49(s29[50],c29[50],andpr32[49],c30[50],s30[49]);


full_add fa30_50(s29[51],c29[51],andpr32[50],c30[51],s30[50]);


full_add fa30_51(s29[52],c29[52],andpr32[51],c30[52],s30[51]);


full_add fa30_52(s29[53],c29[53],andpr32[52],c30[53],s30[52]);


full_add fa30_53(s29[54],c29[54],andpr32[53],c30[54],s30[53]);


full_add fa30_54(s29[55],c29[55],andpr32[54],c30[55],s30[54]);


full_add fa30_55(s29[56],c29[56],andpr32[55],c30[56],s30[55]);


full_add fa30_56(s29[57],c29[57],andpr32[56],c30[57],s30[56]);


full_add fa30_57(s29[58],c29[58],andpr32[57],c30[58],s30[57]);


full_add fa30_58(s29[59],c29[59],andpr32[58],c30[59],s30[58]);


full_add fa30_59(s29[60],c29[60],andpr32[59],c30[60],s30[59]);


full_add fa30_60(s29[61],c29[61],andpr32[60],c30[61],s30[60]);


full_add fa30_61(s29[62],c29[62],andpr32[61],c30[62],s30[61]);


full_add fa30_62(si[30],c29[63],andpr32[62],c30[63],s30[62]);



half_adder ha31(s30[0],c30[0],c31[0],p[31]);


full_add fa31_0(s30[1],c30[1],andpr33[0],c31[1],s31[0]);


full_add fa31_1(s30[2],c30[2],andpr33[1],c31[2],s31[1]);


full_add fa31_2(s30[3],c30[3],andpr33[2],c31[3],s31[2]);


full_add fa31_3(s30[4],c30[4],andpr33[3],c31[4],s31[3]);


full_add fa31_4(s30[5],c30[5],andpr33[4],c31[5],s31[4]);


full_add fa31_5(s30[6],c30[6],andpr33[5],c31[6],s31[5]);


full_add fa31_6(s30[7],c30[7],andpr33[6],c31[7],s31[6]);


full_add fa31_7(s30[8],c30[8],andpr33[7],c31[8],s31[7]);


full_add fa31_8(s30[9],c30[9],andpr33[8],c31[9],s31[8]);


full_add fa31_9(s30[10],c30[10],andpr33[9],c31[10],s31[9]);


full_add fa31_10(s30[11],c30[11],andpr33[10],c31[11],s31[10]);


full_add fa31_11(s30[12],c30[12],andpr33[11],c31[12],s31[11]);


full_add fa31_12(s30[13],c30[13],andpr33[12],c31[13],s31[12]);


full_add fa31_13(s30[14],c30[14],andpr33[13],c31[14],s31[13]);


full_add fa31_14(s30[15],c30[15],andpr33[14],c31[15],s31[14]);


full_add fa31_15(s30[16],c30[16],andpr33[15],c31[16],s31[15]);


full_add fa31_16(s30[17],c30[17],andpr33[16],c31[17],s31[16]);


full_add fa31_17(s30[18],c30[18],andpr33[17],c31[18],s31[17]);


full_add fa31_18(s30[19],c30[19],andpr33[18],c31[19],s31[18]);


full_add fa31_19(s30[20],c30[20],andpr33[19],c31[20],s31[19]);


full_add fa31_20(s30[21],c30[21],andpr33[20],c31[21],s31[20]);


full_add fa31_21(s30[22],c30[22],andpr33[21],c31[22],s31[21]);


full_add fa31_22(s30[23],c30[23],andpr33[22],c31[23],s31[22]);


full_add fa31_23(s30[24],c30[24],andpr33[23],c31[24],s31[23]);


full_add fa31_24(s30[25],c30[25],andpr33[24],c31[25],s31[24]);


full_add fa31_25(s30[26],c30[26],andpr33[25],c31[26],s31[25]);


full_add fa31_26(s30[27],c30[27],andpr33[26],c31[27],s31[26]);


full_add fa31_27(s30[28],c30[28],andpr33[27],c31[28],s31[27]);


full_add fa31_28(s30[29],c30[29],andpr33[28],c31[29],s31[28]);


full_add fa31_29(s30[30],c30[30],andpr33[29],c31[30],s31[29]);


full_add fa31_30(s30[31],c30[31],andpr33[30],c31[31],s31[30]);


full_add fa31_31(s30[32],c30[32],andpr33[31],c31[32],s31[31]);


full_add fa31_32(s30[33],c30[33],andpr33[32],c31[33],s31[32]);


full_add fa31_33(s30[34],c30[34],andpr33[33],c31[34],s31[33]);


full_add fa31_34(s30[35],c30[35],andpr33[34],c31[35],s31[34]);


full_add fa31_35(s30[36],c30[36],andpr33[35],c31[36],s31[35]);


full_add fa31_36(s30[37],c30[37],andpr33[36],c31[37],s31[36]);


full_add fa31_37(s30[38],c30[38],andpr33[37],c31[38],s31[37]);


full_add fa31_38(s30[39],c30[39],andpr33[38],c31[39],s31[38]);


full_add fa31_39(s30[40],c30[40],andpr33[39],c31[40],s31[39]);


full_add fa31_40(s30[41],c30[41],andpr33[40],c31[41],s31[40]);


full_add fa31_41(s30[42],c30[42],andpr33[41],c31[42],s31[41]);


full_add fa31_42(s30[43],c30[43],andpr33[42],c31[43],s31[42]);


full_add fa31_43(s30[44],c30[44],andpr33[43],c31[44],s31[43]);


full_add fa31_44(s30[45],c30[45],andpr33[44],c31[45],s31[44]);


full_add fa31_45(s30[46],c30[46],andpr33[45],c31[46],s31[45]);


full_add fa31_46(s30[47],c30[47],andpr33[46],c31[47],s31[46]);


full_add fa31_47(s30[48],c30[48],andpr33[47],c31[48],s31[47]);


full_add fa31_48(s30[49],c30[49],andpr33[48],c31[49],s31[48]);


full_add fa31_49(s30[50],c30[50],andpr33[49],c31[50],s31[49]);


full_add fa31_50(s30[51],c30[51],andpr33[50],c31[51],s31[50]);


full_add fa31_51(s30[52],c30[52],andpr33[51],c31[52],s31[51]);


full_add fa31_52(s30[53],c30[53],andpr33[52],c31[53],s31[52]);


full_add fa31_53(s30[54],c30[54],andpr33[53],c31[54],s31[53]);


full_add fa31_54(s30[55],c30[55],andpr33[54],c31[55],s31[54]);


full_add fa31_55(s30[56],c30[56],andpr33[55],c31[56],s31[55]);


full_add fa31_56(s30[57],c30[57],andpr33[56],c31[57],s31[56]);


full_add fa31_57(s30[58],c30[58],andpr33[57],c31[58],s31[57]);


full_add fa31_58(s30[59],c30[59],andpr33[58],c31[59],s31[58]);


full_add fa31_59(s30[60],c30[60],andpr33[59],c31[60],s31[59]);


full_add fa31_60(s30[61],c30[61],andpr33[60],c31[61],s31[60]);


full_add fa31_61(s30[62],c30[62],andpr33[61],c31[62],s31[61]);


full_add fa31_62(si[31],c30[63],andpr33[62],c31[63],s31[62]);



half_adder ha32(s31[0],c31[0],c32[0],p[32]);


full_add fa32_0(s31[1],c31[1],andpr34[0],c32[1],s32[0]);


full_add fa32_1(s31[2],c31[2],andpr34[1],c32[2],s32[1]);


full_add fa32_2(s31[3],c31[3],andpr34[2],c32[3],s32[2]);


full_add fa32_3(s31[4],c31[4],andpr34[3],c32[4],s32[3]);


full_add fa32_4(s31[5],c31[5],andpr34[4],c32[5],s32[4]);


full_add fa32_5(s31[6],c31[6],andpr34[5],c32[6],s32[5]);


full_add fa32_6(s31[7],c31[7],andpr34[6],c32[7],s32[6]);


full_add fa32_7(s31[8],c31[8],andpr34[7],c32[8],s32[7]);


full_add fa32_8(s31[9],c31[9],andpr34[8],c32[9],s32[8]);


full_add fa32_9(s31[10],c31[10],andpr34[9],c32[10],s32[9]);


full_add fa32_10(s31[11],c31[11],andpr34[10],c32[11],s32[10]);


full_add fa32_11(s31[12],c31[12],andpr34[11],c32[12],s32[11]);


full_add fa32_12(s31[13],c31[13],andpr34[12],c32[13],s32[12]);


full_add fa32_13(s31[14],c31[14],andpr34[13],c32[14],s32[13]);


full_add fa32_14(s31[15],c31[15],andpr34[14],c32[15],s32[14]);


full_add fa32_15(s31[16],c31[16],andpr34[15],c32[16],s32[15]);


full_add fa32_16(s31[17],c31[17],andpr34[16],c32[17],s32[16]);


full_add fa32_17(s31[18],c31[18],andpr34[17],c32[18],s32[17]);


full_add fa32_18(s31[19],c31[19],andpr34[18],c32[19],s32[18]);


full_add fa32_19(s31[20],c31[20],andpr34[19],c32[20],s32[19]);


full_add fa32_20(s31[21],c31[21],andpr34[20],c32[21],s32[20]);


full_add fa32_21(s31[22],c31[22],andpr34[21],c32[22],s32[21]);


full_add fa32_22(s31[23],c31[23],andpr34[22],c32[23],s32[22]);


full_add fa32_23(s31[24],c31[24],andpr34[23],c32[24],s32[23]);


full_add fa32_24(s31[25],c31[25],andpr34[24],c32[25],s32[24]);


full_add fa32_25(s31[26],c31[26],andpr34[25],c32[26],s32[25]);


full_add fa32_26(s31[27],c31[27],andpr34[26],c32[27],s32[26]);


full_add fa32_27(s31[28],c31[28],andpr34[27],c32[28],s32[27]);


full_add fa32_28(s31[29],c31[29],andpr34[28],c32[29],s32[28]);


full_add fa32_29(s31[30],c31[30],andpr34[29],c32[30],s32[29]);


full_add fa32_30(s31[31],c31[31],andpr34[30],c32[31],s32[30]);


full_add fa32_31(s31[32],c31[32],andpr34[31],c32[32],s32[31]);


full_add fa32_32(s31[33],c31[33],andpr34[32],c32[33],s32[32]);


full_add fa32_33(s31[34],c31[34],andpr34[33],c32[34],s32[33]);


full_add fa32_34(s31[35],c31[35],andpr34[34],c32[35],s32[34]);


full_add fa32_35(s31[36],c31[36],andpr34[35],c32[36],s32[35]);


full_add fa32_36(s31[37],c31[37],andpr34[36],c32[37],s32[36]);


full_add fa32_37(s31[38],c31[38],andpr34[37],c32[38],s32[37]);


full_add fa32_38(s31[39],c31[39],andpr34[38],c32[39],s32[38]);


full_add fa32_39(s31[40],c31[40],andpr34[39],c32[40],s32[39]);


full_add fa32_40(s31[41],c31[41],andpr34[40],c32[41],s32[40]);


full_add fa32_41(s31[42],c31[42],andpr34[41],c32[42],s32[41]);


full_add fa32_42(s31[43],c31[43],andpr34[42],c32[43],s32[42]);


full_add fa32_43(s31[44],c31[44],andpr34[43],c32[44],s32[43]);


full_add fa32_44(s31[45],c31[45],andpr34[44],c32[45],s32[44]);


full_add fa32_45(s31[46],c31[46],andpr34[45],c32[46],s32[45]);


full_add fa32_46(s31[47],c31[47],andpr34[46],c32[47],s32[46]);


full_add fa32_47(s31[48],c31[48],andpr34[47],c32[48],s32[47]);


full_add fa32_48(s31[49],c31[49],andpr34[48],c32[49],s32[48]);


full_add fa32_49(s31[50],c31[50],andpr34[49],c32[50],s32[49]);


full_add fa32_50(s31[51],c31[51],andpr34[50],c32[51],s32[50]);


full_add fa32_51(s31[52],c31[52],andpr34[51],c32[52],s32[51]);


full_add fa32_52(s31[53],c31[53],andpr34[52],c32[53],s32[52]);


full_add fa32_53(s31[54],c31[54],andpr34[53],c32[54],s32[53]);


full_add fa32_54(s31[55],c31[55],andpr34[54],c32[55],s32[54]);


full_add fa32_55(s31[56],c31[56],andpr34[55],c32[56],s32[55]);


full_add fa32_56(s31[57],c31[57],andpr34[56],c32[57],s32[56]);


full_add fa32_57(s31[58],c31[58],andpr34[57],c32[58],s32[57]);


full_add fa32_58(s31[59],c31[59],andpr34[58],c32[59],s32[58]);


full_add fa32_59(s31[60],c31[60],andpr34[59],c32[60],s32[59]);


full_add fa32_60(s31[61],c31[61],andpr34[60],c32[61],s32[60]);


full_add fa32_61(s31[62],c31[62],andpr34[61],c32[62],s32[61]);


full_add fa32_62(si[32],c31[63],andpr34[62],c32[63],s32[62]);



half_adder ha33(s32[0],c32[0],c33[0],p[33]);


full_add fa33_0(s32[1],c32[1],andpr35[0],c33[1],s33[0]);


full_add fa33_1(s32[2],c32[2],andpr35[1],c33[2],s33[1]);


full_add fa33_2(s32[3],c32[3],andpr35[2],c33[3],s33[2]);


full_add fa33_3(s32[4],c32[4],andpr35[3],c33[4],s33[3]);


full_add fa33_4(s32[5],c32[5],andpr35[4],c33[5],s33[4]);


full_add fa33_5(s32[6],c32[6],andpr35[5],c33[6],s33[5]);


full_add fa33_6(s32[7],c32[7],andpr35[6],c33[7],s33[6]);


full_add fa33_7(s32[8],c32[8],andpr35[7],c33[8],s33[7]);


full_add fa33_8(s32[9],c32[9],andpr35[8],c33[9],s33[8]);


full_add fa33_9(s32[10],c32[10],andpr35[9],c33[10],s33[9]);


full_add fa33_10(s32[11],c32[11],andpr35[10],c33[11],s33[10]);


full_add fa33_11(s32[12],c32[12],andpr35[11],c33[12],s33[11]);


full_add fa33_12(s32[13],c32[13],andpr35[12],c33[13],s33[12]);


full_add fa33_13(s32[14],c32[14],andpr35[13],c33[14],s33[13]);


full_add fa33_14(s32[15],c32[15],andpr35[14],c33[15],s33[14]);


full_add fa33_15(s32[16],c32[16],andpr35[15],c33[16],s33[15]);


full_add fa33_16(s32[17],c32[17],andpr35[16],c33[17],s33[16]);


full_add fa33_17(s32[18],c32[18],andpr35[17],c33[18],s33[17]);


full_add fa33_18(s32[19],c32[19],andpr35[18],c33[19],s33[18]);


full_add fa33_19(s32[20],c32[20],andpr35[19],c33[20],s33[19]);


full_add fa33_20(s32[21],c32[21],andpr35[20],c33[21],s33[20]);


full_add fa33_21(s32[22],c32[22],andpr35[21],c33[22],s33[21]);


full_add fa33_22(s32[23],c32[23],andpr35[22],c33[23],s33[22]);


full_add fa33_23(s32[24],c32[24],andpr35[23],c33[24],s33[23]);


full_add fa33_24(s32[25],c32[25],andpr35[24],c33[25],s33[24]);


full_add fa33_25(s32[26],c32[26],andpr35[25],c33[26],s33[25]);


full_add fa33_26(s32[27],c32[27],andpr35[26],c33[27],s33[26]);


full_add fa33_27(s32[28],c32[28],andpr35[27],c33[28],s33[27]);


full_add fa33_28(s32[29],c32[29],andpr35[28],c33[29],s33[28]);


full_add fa33_29(s32[30],c32[30],andpr35[29],c33[30],s33[29]);


full_add fa33_30(s32[31],c32[31],andpr35[30],c33[31],s33[30]);


full_add fa33_31(s32[32],c32[32],andpr35[31],c33[32],s33[31]);


full_add fa33_32(s32[33],c32[33],andpr35[32],c33[33],s33[32]);


full_add fa33_33(s32[34],c32[34],andpr35[33],c33[34],s33[33]);


full_add fa33_34(s32[35],c32[35],andpr35[34],c33[35],s33[34]);


full_add fa33_35(s32[36],c32[36],andpr35[35],c33[36],s33[35]);


full_add fa33_36(s32[37],c32[37],andpr35[36],c33[37],s33[36]);


full_add fa33_37(s32[38],c32[38],andpr35[37],c33[38],s33[37]);


full_add fa33_38(s32[39],c32[39],andpr35[38],c33[39],s33[38]);


full_add fa33_39(s32[40],c32[40],andpr35[39],c33[40],s33[39]);


full_add fa33_40(s32[41],c32[41],andpr35[40],c33[41],s33[40]);


full_add fa33_41(s32[42],c32[42],andpr35[41],c33[42],s33[41]);


full_add fa33_42(s32[43],c32[43],andpr35[42],c33[43],s33[42]);


full_add fa33_43(s32[44],c32[44],andpr35[43],c33[44],s33[43]);


full_add fa33_44(s32[45],c32[45],andpr35[44],c33[45],s33[44]);


full_add fa33_45(s32[46],c32[46],andpr35[45],c33[46],s33[45]);


full_add fa33_46(s32[47],c32[47],andpr35[46],c33[47],s33[46]);


full_add fa33_47(s32[48],c32[48],andpr35[47],c33[48],s33[47]);


full_add fa33_48(s32[49],c32[49],andpr35[48],c33[49],s33[48]);


full_add fa33_49(s32[50],c32[50],andpr35[49],c33[50],s33[49]);


full_add fa33_50(s32[51],c32[51],andpr35[50],c33[51],s33[50]);


full_add fa33_51(s32[52],c32[52],andpr35[51],c33[52],s33[51]);


full_add fa33_52(s32[53],c32[53],andpr35[52],c33[53],s33[52]);


full_add fa33_53(s32[54],c32[54],andpr35[53],c33[54],s33[53]);


full_add fa33_54(s32[55],c32[55],andpr35[54],c33[55],s33[54]);


full_add fa33_55(s32[56],c32[56],andpr35[55],c33[56],s33[55]);


full_add fa33_56(s32[57],c32[57],andpr35[56],c33[57],s33[56]);


full_add fa33_57(s32[58],c32[58],andpr35[57],c33[58],s33[57]);


full_add fa33_58(s32[59],c32[59],andpr35[58],c33[59],s33[58]);


full_add fa33_59(s32[60],c32[60],andpr35[59],c33[60],s33[59]);


full_add fa33_60(s32[61],c32[61],andpr35[60],c33[61],s33[60]);


full_add fa33_61(s32[62],c32[62],andpr35[61],c33[62],s33[61]);


full_add fa33_62(si[33],c32[63],andpr35[62],c33[63],s33[62]);



half_adder ha34(s33[0],c33[0],c34[0],p[34]);


full_add fa34_0(s33[1],c33[1],andpr36[0],c34[1],s34[0]);


full_add fa34_1(s33[2],c33[2],andpr36[1],c34[2],s34[1]);


full_add fa34_2(s33[3],c33[3],andpr36[2],c34[3],s34[2]);


full_add fa34_3(s33[4],c33[4],andpr36[3],c34[4],s34[3]);


full_add fa34_4(s33[5],c33[5],andpr36[4],c34[5],s34[4]);


full_add fa34_5(s33[6],c33[6],andpr36[5],c34[6],s34[5]);


full_add fa34_6(s33[7],c33[7],andpr36[6],c34[7],s34[6]);


full_add fa34_7(s33[8],c33[8],andpr36[7],c34[8],s34[7]);


full_add fa34_8(s33[9],c33[9],andpr36[8],c34[9],s34[8]);


full_add fa34_9(s33[10],c33[10],andpr36[9],c34[10],s34[9]);


full_add fa34_10(s33[11],c33[11],andpr36[10],c34[11],s34[10]);


full_add fa34_11(s33[12],c33[12],andpr36[11],c34[12],s34[11]);


full_add fa34_12(s33[13],c33[13],andpr36[12],c34[13],s34[12]);


full_add fa34_13(s33[14],c33[14],andpr36[13],c34[14],s34[13]);


full_add fa34_14(s33[15],c33[15],andpr36[14],c34[15],s34[14]);


full_add fa34_15(s33[16],c33[16],andpr36[15],c34[16],s34[15]);


full_add fa34_16(s33[17],c33[17],andpr36[16],c34[17],s34[16]);


full_add fa34_17(s33[18],c33[18],andpr36[17],c34[18],s34[17]);


full_add fa34_18(s33[19],c33[19],andpr36[18],c34[19],s34[18]);


full_add fa34_19(s33[20],c33[20],andpr36[19],c34[20],s34[19]);


full_add fa34_20(s33[21],c33[21],andpr36[20],c34[21],s34[20]);


full_add fa34_21(s33[22],c33[22],andpr36[21],c34[22],s34[21]);


full_add fa34_22(s33[23],c33[23],andpr36[22],c34[23],s34[22]);


full_add fa34_23(s33[24],c33[24],andpr36[23],c34[24],s34[23]);


full_add fa34_24(s33[25],c33[25],andpr36[24],c34[25],s34[24]);


full_add fa34_25(s33[26],c33[26],andpr36[25],c34[26],s34[25]);


full_add fa34_26(s33[27],c33[27],andpr36[26],c34[27],s34[26]);


full_add fa34_27(s33[28],c33[28],andpr36[27],c34[28],s34[27]);


full_add fa34_28(s33[29],c33[29],andpr36[28],c34[29],s34[28]);


full_add fa34_29(s33[30],c33[30],andpr36[29],c34[30],s34[29]);


full_add fa34_30(s33[31],c33[31],andpr36[30],c34[31],s34[30]);


full_add fa34_31(s33[32],c33[32],andpr36[31],c34[32],s34[31]);


full_add fa34_32(s33[33],c33[33],andpr36[32],c34[33],s34[32]);


full_add fa34_33(s33[34],c33[34],andpr36[33],c34[34],s34[33]);


full_add fa34_34(s33[35],c33[35],andpr36[34],c34[35],s34[34]);


full_add fa34_35(s33[36],c33[36],andpr36[35],c34[36],s34[35]);


full_add fa34_36(s33[37],c33[37],andpr36[36],c34[37],s34[36]);


full_add fa34_37(s33[38],c33[38],andpr36[37],c34[38],s34[37]);


full_add fa34_38(s33[39],c33[39],andpr36[38],c34[39],s34[38]);


full_add fa34_39(s33[40],c33[40],andpr36[39],c34[40],s34[39]);


full_add fa34_40(s33[41],c33[41],andpr36[40],c34[41],s34[40]);


full_add fa34_41(s33[42],c33[42],andpr36[41],c34[42],s34[41]);


full_add fa34_42(s33[43],c33[43],andpr36[42],c34[43],s34[42]);


full_add fa34_43(s33[44],c33[44],andpr36[43],c34[44],s34[43]);


full_add fa34_44(s33[45],c33[45],andpr36[44],c34[45],s34[44]);


full_add fa34_45(s33[46],c33[46],andpr36[45],c34[46],s34[45]);


full_add fa34_46(s33[47],c33[47],andpr36[46],c34[47],s34[46]);


full_add fa34_47(s33[48],c33[48],andpr36[47],c34[48],s34[47]);


full_add fa34_48(s33[49],c33[49],andpr36[48],c34[49],s34[48]);


full_add fa34_49(s33[50],c33[50],andpr36[49],c34[50],s34[49]);


full_add fa34_50(s33[51],c33[51],andpr36[50],c34[51],s34[50]);


full_add fa34_51(s33[52],c33[52],andpr36[51],c34[52],s34[51]);


full_add fa34_52(s33[53],c33[53],andpr36[52],c34[53],s34[52]);


full_add fa34_53(s33[54],c33[54],andpr36[53],c34[54],s34[53]);


full_add fa34_54(s33[55],c33[55],andpr36[54],c34[55],s34[54]);


full_add fa34_55(s33[56],c33[56],andpr36[55],c34[56],s34[55]);


full_add fa34_56(s33[57],c33[57],andpr36[56],c34[57],s34[56]);


full_add fa34_57(s33[58],c33[58],andpr36[57],c34[58],s34[57]);


full_add fa34_58(s33[59],c33[59],andpr36[58],c34[59],s34[58]);


full_add fa34_59(s33[60],c33[60],andpr36[59],c34[60],s34[59]);


full_add fa34_60(s33[61],c33[61],andpr36[60],c34[61],s34[60]);


full_add fa34_61(s33[62],c33[62],andpr36[61],c34[62],s34[61]);


full_add fa34_62(si[34],c33[63],andpr36[62],c34[63],s34[62]);



half_adder ha35(s34[0],c34[0],c35[0],p[35]);


full_add fa35_0(s34[1],c34[1],andpr37[0],c35[1],s35[0]);


full_add fa35_1(s34[2],c34[2],andpr37[1],c35[2],s35[1]);


full_add fa35_2(s34[3],c34[3],andpr37[2],c35[3],s35[2]);


full_add fa35_3(s34[4],c34[4],andpr37[3],c35[4],s35[3]);


full_add fa35_4(s34[5],c34[5],andpr37[4],c35[5],s35[4]);


full_add fa35_5(s34[6],c34[6],andpr37[5],c35[6],s35[5]);


full_add fa35_6(s34[7],c34[7],andpr37[6],c35[7],s35[6]);


full_add fa35_7(s34[8],c34[8],andpr37[7],c35[8],s35[7]);


full_add fa35_8(s34[9],c34[9],andpr37[8],c35[9],s35[8]);


full_add fa35_9(s34[10],c34[10],andpr37[9],c35[10],s35[9]);


full_add fa35_10(s34[11],c34[11],andpr37[10],c35[11],s35[10]);


full_add fa35_11(s34[12],c34[12],andpr37[11],c35[12],s35[11]);


full_add fa35_12(s34[13],c34[13],andpr37[12],c35[13],s35[12]);


full_add fa35_13(s34[14],c34[14],andpr37[13],c35[14],s35[13]);


full_add fa35_14(s34[15],c34[15],andpr37[14],c35[15],s35[14]);


full_add fa35_15(s34[16],c34[16],andpr37[15],c35[16],s35[15]);


full_add fa35_16(s34[17],c34[17],andpr37[16],c35[17],s35[16]);


full_add fa35_17(s34[18],c34[18],andpr37[17],c35[18],s35[17]);


full_add fa35_18(s34[19],c34[19],andpr37[18],c35[19],s35[18]);


full_add fa35_19(s34[20],c34[20],andpr37[19],c35[20],s35[19]);


full_add fa35_20(s34[21],c34[21],andpr37[20],c35[21],s35[20]);


full_add fa35_21(s34[22],c34[22],andpr37[21],c35[22],s35[21]);


full_add fa35_22(s34[23],c34[23],andpr37[22],c35[23],s35[22]);


full_add fa35_23(s34[24],c34[24],andpr37[23],c35[24],s35[23]);


full_add fa35_24(s34[25],c34[25],andpr37[24],c35[25],s35[24]);


full_add fa35_25(s34[26],c34[26],andpr37[25],c35[26],s35[25]);


full_add fa35_26(s34[27],c34[27],andpr37[26],c35[27],s35[26]);


full_add fa35_27(s34[28],c34[28],andpr37[27],c35[28],s35[27]);


full_add fa35_28(s34[29],c34[29],andpr37[28],c35[29],s35[28]);


full_add fa35_29(s34[30],c34[30],andpr37[29],c35[30],s35[29]);


full_add fa35_30(s34[31],c34[31],andpr37[30],c35[31],s35[30]);


full_add fa35_31(s34[32],c34[32],andpr37[31],c35[32],s35[31]);


full_add fa35_32(s34[33],c34[33],andpr37[32],c35[33],s35[32]);


full_add fa35_33(s34[34],c34[34],andpr37[33],c35[34],s35[33]);


full_add fa35_34(s34[35],c34[35],andpr37[34],c35[35],s35[34]);


full_add fa35_35(s34[36],c34[36],andpr37[35],c35[36],s35[35]);


full_add fa35_36(s34[37],c34[37],andpr37[36],c35[37],s35[36]);


full_add fa35_37(s34[38],c34[38],andpr37[37],c35[38],s35[37]);


full_add fa35_38(s34[39],c34[39],andpr37[38],c35[39],s35[38]);


full_add fa35_39(s34[40],c34[40],andpr37[39],c35[40],s35[39]);


full_add fa35_40(s34[41],c34[41],andpr37[40],c35[41],s35[40]);


full_add fa35_41(s34[42],c34[42],andpr37[41],c35[42],s35[41]);


full_add fa35_42(s34[43],c34[43],andpr37[42],c35[43],s35[42]);


full_add fa35_43(s34[44],c34[44],andpr37[43],c35[44],s35[43]);


full_add fa35_44(s34[45],c34[45],andpr37[44],c35[45],s35[44]);


full_add fa35_45(s34[46],c34[46],andpr37[45],c35[46],s35[45]);


full_add fa35_46(s34[47],c34[47],andpr37[46],c35[47],s35[46]);


full_add fa35_47(s34[48],c34[48],andpr37[47],c35[48],s35[47]);


full_add fa35_48(s34[49],c34[49],andpr37[48],c35[49],s35[48]);


full_add fa35_49(s34[50],c34[50],andpr37[49],c35[50],s35[49]);


full_add fa35_50(s34[51],c34[51],andpr37[50],c35[51],s35[50]);


full_add fa35_51(s34[52],c34[52],andpr37[51],c35[52],s35[51]);


full_add fa35_52(s34[53],c34[53],andpr37[52],c35[53],s35[52]);


full_add fa35_53(s34[54],c34[54],andpr37[53],c35[54],s35[53]);


full_add fa35_54(s34[55],c34[55],andpr37[54],c35[55],s35[54]);


full_add fa35_55(s34[56],c34[56],andpr37[55],c35[56],s35[55]);


full_add fa35_56(s34[57],c34[57],andpr37[56],c35[57],s35[56]);


full_add fa35_57(s34[58],c34[58],andpr37[57],c35[58],s35[57]);


full_add fa35_58(s34[59],c34[59],andpr37[58],c35[59],s35[58]);


full_add fa35_59(s34[60],c34[60],andpr37[59],c35[60],s35[59]);


full_add fa35_60(s34[61],c34[61],andpr37[60],c35[61],s35[60]);


full_add fa35_61(s34[62],c34[62],andpr37[61],c35[62],s35[61]);


full_add fa35_62(si[35],c34[63],andpr37[62],c35[63],s35[62]);



half_adder ha36(s35[0],c35[0],c36[0],p[36]);


full_add fa36_0(s35[1],c35[1],andpr38[0],c36[1],s36[0]);


full_add fa36_1(s35[2],c35[2],andpr38[1],c36[2],s36[1]);


full_add fa36_2(s35[3],c35[3],andpr38[2],c36[3],s36[2]);


full_add fa36_3(s35[4],c35[4],andpr38[3],c36[4],s36[3]);


full_add fa36_4(s35[5],c35[5],andpr38[4],c36[5],s36[4]);


full_add fa36_5(s35[6],c35[6],andpr38[5],c36[6],s36[5]);


full_add fa36_6(s35[7],c35[7],andpr38[6],c36[7],s36[6]);


full_add fa36_7(s35[8],c35[8],andpr38[7],c36[8],s36[7]);


full_add fa36_8(s35[9],c35[9],andpr38[8],c36[9],s36[8]);


full_add fa36_9(s35[10],c35[10],andpr38[9],c36[10],s36[9]);


full_add fa36_10(s35[11],c35[11],andpr38[10],c36[11],s36[10]);


full_add fa36_11(s35[12],c35[12],andpr38[11],c36[12],s36[11]);


full_add fa36_12(s35[13],c35[13],andpr38[12],c36[13],s36[12]);


full_add fa36_13(s35[14],c35[14],andpr38[13],c36[14],s36[13]);


full_add fa36_14(s35[15],c35[15],andpr38[14],c36[15],s36[14]);


full_add fa36_15(s35[16],c35[16],andpr38[15],c36[16],s36[15]);


full_add fa36_16(s35[17],c35[17],andpr38[16],c36[17],s36[16]);


full_add fa36_17(s35[18],c35[18],andpr38[17],c36[18],s36[17]);


full_add fa36_18(s35[19],c35[19],andpr38[18],c36[19],s36[18]);


full_add fa36_19(s35[20],c35[20],andpr38[19],c36[20],s36[19]);


full_add fa36_20(s35[21],c35[21],andpr38[20],c36[21],s36[20]);


full_add fa36_21(s35[22],c35[22],andpr38[21],c36[22],s36[21]);


full_add fa36_22(s35[23],c35[23],andpr38[22],c36[23],s36[22]);


full_add fa36_23(s35[24],c35[24],andpr38[23],c36[24],s36[23]);


full_add fa36_24(s35[25],c35[25],andpr38[24],c36[25],s36[24]);


full_add fa36_25(s35[26],c35[26],andpr38[25],c36[26],s36[25]);


full_add fa36_26(s35[27],c35[27],andpr38[26],c36[27],s36[26]);


full_add fa36_27(s35[28],c35[28],andpr38[27],c36[28],s36[27]);


full_add fa36_28(s35[29],c35[29],andpr38[28],c36[29],s36[28]);


full_add fa36_29(s35[30],c35[30],andpr38[29],c36[30],s36[29]);


full_add fa36_30(s35[31],c35[31],andpr38[30],c36[31],s36[30]);


full_add fa36_31(s35[32],c35[32],andpr38[31],c36[32],s36[31]);


full_add fa36_32(s35[33],c35[33],andpr38[32],c36[33],s36[32]);


full_add fa36_33(s35[34],c35[34],andpr38[33],c36[34],s36[33]);


full_add fa36_34(s35[35],c35[35],andpr38[34],c36[35],s36[34]);


full_add fa36_35(s35[36],c35[36],andpr38[35],c36[36],s36[35]);


full_add fa36_36(s35[37],c35[37],andpr38[36],c36[37],s36[36]);


full_add fa36_37(s35[38],c35[38],andpr38[37],c36[38],s36[37]);


full_add fa36_38(s35[39],c35[39],andpr38[38],c36[39],s36[38]);


full_add fa36_39(s35[40],c35[40],andpr38[39],c36[40],s36[39]);


full_add fa36_40(s35[41],c35[41],andpr38[40],c36[41],s36[40]);


full_add fa36_41(s35[42],c35[42],andpr38[41],c36[42],s36[41]);


full_add fa36_42(s35[43],c35[43],andpr38[42],c36[43],s36[42]);


full_add fa36_43(s35[44],c35[44],andpr38[43],c36[44],s36[43]);


full_add fa36_44(s35[45],c35[45],andpr38[44],c36[45],s36[44]);


full_add fa36_45(s35[46],c35[46],andpr38[45],c36[46],s36[45]);


full_add fa36_46(s35[47],c35[47],andpr38[46],c36[47],s36[46]);


full_add fa36_47(s35[48],c35[48],andpr38[47],c36[48],s36[47]);


full_add fa36_48(s35[49],c35[49],andpr38[48],c36[49],s36[48]);


full_add fa36_49(s35[50],c35[50],andpr38[49],c36[50],s36[49]);


full_add fa36_50(s35[51],c35[51],andpr38[50],c36[51],s36[50]);


full_add fa36_51(s35[52],c35[52],andpr38[51],c36[52],s36[51]);


full_add fa36_52(s35[53],c35[53],andpr38[52],c36[53],s36[52]);


full_add fa36_53(s35[54],c35[54],andpr38[53],c36[54],s36[53]);


full_add fa36_54(s35[55],c35[55],andpr38[54],c36[55],s36[54]);


full_add fa36_55(s35[56],c35[56],andpr38[55],c36[56],s36[55]);


full_add fa36_56(s35[57],c35[57],andpr38[56],c36[57],s36[56]);


full_add fa36_57(s35[58],c35[58],andpr38[57],c36[58],s36[57]);


full_add fa36_58(s35[59],c35[59],andpr38[58],c36[59],s36[58]);


full_add fa36_59(s35[60],c35[60],andpr38[59],c36[60],s36[59]);


full_add fa36_60(s35[61],c35[61],andpr38[60],c36[61],s36[60]);


full_add fa36_61(s35[62],c35[62],andpr38[61],c36[62],s36[61]);


full_add fa36_62(si[36],c35[63],andpr38[62],c36[63],s36[62]);



half_adder ha37(s36[0],c36[0],c37[0],p[37]);


full_add fa37_0(s36[1],c36[1],andpr39[0],c37[1],s37[0]);


full_add fa37_1(s36[2],c36[2],andpr39[1],c37[2],s37[1]);


full_add fa37_2(s36[3],c36[3],andpr39[2],c37[3],s37[2]);


full_add fa37_3(s36[4],c36[4],andpr39[3],c37[4],s37[3]);


full_add fa37_4(s36[5],c36[5],andpr39[4],c37[5],s37[4]);


full_add fa37_5(s36[6],c36[6],andpr39[5],c37[6],s37[5]);


full_add fa37_6(s36[7],c36[7],andpr39[6],c37[7],s37[6]);


full_add fa37_7(s36[8],c36[8],andpr39[7],c37[8],s37[7]);


full_add fa37_8(s36[9],c36[9],andpr39[8],c37[9],s37[8]);


full_add fa37_9(s36[10],c36[10],andpr39[9],c37[10],s37[9]);


full_add fa37_10(s36[11],c36[11],andpr39[10],c37[11],s37[10]);


full_add fa37_11(s36[12],c36[12],andpr39[11],c37[12],s37[11]);


full_add fa37_12(s36[13],c36[13],andpr39[12],c37[13],s37[12]);


full_add fa37_13(s36[14],c36[14],andpr39[13],c37[14],s37[13]);


full_add fa37_14(s36[15],c36[15],andpr39[14],c37[15],s37[14]);


full_add fa37_15(s36[16],c36[16],andpr39[15],c37[16],s37[15]);


full_add fa37_16(s36[17],c36[17],andpr39[16],c37[17],s37[16]);


full_add fa37_17(s36[18],c36[18],andpr39[17],c37[18],s37[17]);


full_add fa37_18(s36[19],c36[19],andpr39[18],c37[19],s37[18]);


full_add fa37_19(s36[20],c36[20],andpr39[19],c37[20],s37[19]);


full_add fa37_20(s36[21],c36[21],andpr39[20],c37[21],s37[20]);


full_add fa37_21(s36[22],c36[22],andpr39[21],c37[22],s37[21]);


full_add fa37_22(s36[23],c36[23],andpr39[22],c37[23],s37[22]);


full_add fa37_23(s36[24],c36[24],andpr39[23],c37[24],s37[23]);


full_add fa37_24(s36[25],c36[25],andpr39[24],c37[25],s37[24]);


full_add fa37_25(s36[26],c36[26],andpr39[25],c37[26],s37[25]);


full_add fa37_26(s36[27],c36[27],andpr39[26],c37[27],s37[26]);


full_add fa37_27(s36[28],c36[28],andpr39[27],c37[28],s37[27]);


full_add fa37_28(s36[29],c36[29],andpr39[28],c37[29],s37[28]);


full_add fa37_29(s36[30],c36[30],andpr39[29],c37[30],s37[29]);


full_add fa37_30(s36[31],c36[31],andpr39[30],c37[31],s37[30]);


full_add fa37_31(s36[32],c36[32],andpr39[31],c37[32],s37[31]);


full_add fa37_32(s36[33],c36[33],andpr39[32],c37[33],s37[32]);


full_add fa37_33(s36[34],c36[34],andpr39[33],c37[34],s37[33]);


full_add fa37_34(s36[35],c36[35],andpr39[34],c37[35],s37[34]);


full_add fa37_35(s36[36],c36[36],andpr39[35],c37[36],s37[35]);


full_add fa37_36(s36[37],c36[37],andpr39[36],c37[37],s37[36]);


full_add fa37_37(s36[38],c36[38],andpr39[37],c37[38],s37[37]);


full_add fa37_38(s36[39],c36[39],andpr39[38],c37[39],s37[38]);


full_add fa37_39(s36[40],c36[40],andpr39[39],c37[40],s37[39]);


full_add fa37_40(s36[41],c36[41],andpr39[40],c37[41],s37[40]);


full_add fa37_41(s36[42],c36[42],andpr39[41],c37[42],s37[41]);


full_add fa37_42(s36[43],c36[43],andpr39[42],c37[43],s37[42]);


full_add fa37_43(s36[44],c36[44],andpr39[43],c37[44],s37[43]);


full_add fa37_44(s36[45],c36[45],andpr39[44],c37[45],s37[44]);


full_add fa37_45(s36[46],c36[46],andpr39[45],c37[46],s37[45]);


full_add fa37_46(s36[47],c36[47],andpr39[46],c37[47],s37[46]);


full_add fa37_47(s36[48],c36[48],andpr39[47],c37[48],s37[47]);


full_add fa37_48(s36[49],c36[49],andpr39[48],c37[49],s37[48]);


full_add fa37_49(s36[50],c36[50],andpr39[49],c37[50],s37[49]);


full_add fa37_50(s36[51],c36[51],andpr39[50],c37[51],s37[50]);


full_add fa37_51(s36[52],c36[52],andpr39[51],c37[52],s37[51]);


full_add fa37_52(s36[53],c36[53],andpr39[52],c37[53],s37[52]);


full_add fa37_53(s36[54],c36[54],andpr39[53],c37[54],s37[53]);


full_add fa37_54(s36[55],c36[55],andpr39[54],c37[55],s37[54]);


full_add fa37_55(s36[56],c36[56],andpr39[55],c37[56],s37[55]);


full_add fa37_56(s36[57],c36[57],andpr39[56],c37[57],s37[56]);


full_add fa37_57(s36[58],c36[58],andpr39[57],c37[58],s37[57]);


full_add fa37_58(s36[59],c36[59],andpr39[58],c37[59],s37[58]);


full_add fa37_59(s36[60],c36[60],andpr39[59],c37[60],s37[59]);


full_add fa37_60(s36[61],c36[61],andpr39[60],c37[61],s37[60]);


full_add fa37_61(s36[62],c36[62],andpr39[61],c37[62],s37[61]);


full_add fa37_62(si[37],c36[63],andpr39[62],c37[63],s37[62]);



half_adder ha38(s37[0],c37[0],c38[0],p[38]);


full_add fa38_0(s37[1],c37[1],andpr40[0],c38[1],s38[0]);


full_add fa38_1(s37[2],c37[2],andpr40[1],c38[2],s38[1]);


full_add fa38_2(s37[3],c37[3],andpr40[2],c38[3],s38[2]);


full_add fa38_3(s37[4],c37[4],andpr40[3],c38[4],s38[3]);


full_add fa38_4(s37[5],c37[5],andpr40[4],c38[5],s38[4]);


full_add fa38_5(s37[6],c37[6],andpr40[5],c38[6],s38[5]);


full_add fa38_6(s37[7],c37[7],andpr40[6],c38[7],s38[6]);


full_add fa38_7(s37[8],c37[8],andpr40[7],c38[8],s38[7]);


full_add fa38_8(s37[9],c37[9],andpr40[8],c38[9],s38[8]);


full_add fa38_9(s37[10],c37[10],andpr40[9],c38[10],s38[9]);


full_add fa38_10(s37[11],c37[11],andpr40[10],c38[11],s38[10]);


full_add fa38_11(s37[12],c37[12],andpr40[11],c38[12],s38[11]);


full_add fa38_12(s37[13],c37[13],andpr40[12],c38[13],s38[12]);


full_add fa38_13(s37[14],c37[14],andpr40[13],c38[14],s38[13]);


full_add fa38_14(s37[15],c37[15],andpr40[14],c38[15],s38[14]);


full_add fa38_15(s37[16],c37[16],andpr40[15],c38[16],s38[15]);


full_add fa38_16(s37[17],c37[17],andpr40[16],c38[17],s38[16]);


full_add fa38_17(s37[18],c37[18],andpr40[17],c38[18],s38[17]);


full_add fa38_18(s37[19],c37[19],andpr40[18],c38[19],s38[18]);


full_add fa38_19(s37[20],c37[20],andpr40[19],c38[20],s38[19]);


full_add fa38_20(s37[21],c37[21],andpr40[20],c38[21],s38[20]);


full_add fa38_21(s37[22],c37[22],andpr40[21],c38[22],s38[21]);


full_add fa38_22(s37[23],c37[23],andpr40[22],c38[23],s38[22]);


full_add fa38_23(s37[24],c37[24],andpr40[23],c38[24],s38[23]);


full_add fa38_24(s37[25],c37[25],andpr40[24],c38[25],s38[24]);


full_add fa38_25(s37[26],c37[26],andpr40[25],c38[26],s38[25]);


full_add fa38_26(s37[27],c37[27],andpr40[26],c38[27],s38[26]);


full_add fa38_27(s37[28],c37[28],andpr40[27],c38[28],s38[27]);


full_add fa38_28(s37[29],c37[29],andpr40[28],c38[29],s38[28]);


full_add fa38_29(s37[30],c37[30],andpr40[29],c38[30],s38[29]);


full_add fa38_30(s37[31],c37[31],andpr40[30],c38[31],s38[30]);


full_add fa38_31(s37[32],c37[32],andpr40[31],c38[32],s38[31]);


full_add fa38_32(s37[33],c37[33],andpr40[32],c38[33],s38[32]);


full_add fa38_33(s37[34],c37[34],andpr40[33],c38[34],s38[33]);


full_add fa38_34(s37[35],c37[35],andpr40[34],c38[35],s38[34]);


full_add fa38_35(s37[36],c37[36],andpr40[35],c38[36],s38[35]);


full_add fa38_36(s37[37],c37[37],andpr40[36],c38[37],s38[36]);


full_add fa38_37(s37[38],c37[38],andpr40[37],c38[38],s38[37]);


full_add fa38_38(s37[39],c37[39],andpr40[38],c38[39],s38[38]);


full_add fa38_39(s37[40],c37[40],andpr40[39],c38[40],s38[39]);


full_add fa38_40(s37[41],c37[41],andpr40[40],c38[41],s38[40]);


full_add fa38_41(s37[42],c37[42],andpr40[41],c38[42],s38[41]);


full_add fa38_42(s37[43],c37[43],andpr40[42],c38[43],s38[42]);


full_add fa38_43(s37[44],c37[44],andpr40[43],c38[44],s38[43]);


full_add fa38_44(s37[45],c37[45],andpr40[44],c38[45],s38[44]);


full_add fa38_45(s37[46],c37[46],andpr40[45],c38[46],s38[45]);


full_add fa38_46(s37[47],c37[47],andpr40[46],c38[47],s38[46]);


full_add fa38_47(s37[48],c37[48],andpr40[47],c38[48],s38[47]);


full_add fa38_48(s37[49],c37[49],andpr40[48],c38[49],s38[48]);


full_add fa38_49(s37[50],c37[50],andpr40[49],c38[50],s38[49]);


full_add fa38_50(s37[51],c37[51],andpr40[50],c38[51],s38[50]);


full_add fa38_51(s37[52],c37[52],andpr40[51],c38[52],s38[51]);


full_add fa38_52(s37[53],c37[53],andpr40[52],c38[53],s38[52]);


full_add fa38_53(s37[54],c37[54],andpr40[53],c38[54],s38[53]);


full_add fa38_54(s37[55],c37[55],andpr40[54],c38[55],s38[54]);


full_add fa38_55(s37[56],c37[56],andpr40[55],c38[56],s38[55]);


full_add fa38_56(s37[57],c37[57],andpr40[56],c38[57],s38[56]);


full_add fa38_57(s37[58],c37[58],andpr40[57],c38[58],s38[57]);


full_add fa38_58(s37[59],c37[59],andpr40[58],c38[59],s38[58]);


full_add fa38_59(s37[60],c37[60],andpr40[59],c38[60],s38[59]);


full_add fa38_60(s37[61],c37[61],andpr40[60],c38[61],s38[60]);


full_add fa38_61(s37[62],c37[62],andpr40[61],c38[62],s38[61]);


full_add fa38_62(si[38],c37[63],andpr40[62],c38[63],s38[62]);



half_adder ha39(s38[0],c38[0],c39[0],p[39]);


full_add fa39_0(s38[1],c38[1],andpr41[0],c39[1],s39[0]);


full_add fa39_1(s38[2],c38[2],andpr41[1],c39[2],s39[1]);


full_add fa39_2(s38[3],c38[3],andpr41[2],c39[3],s39[2]);


full_add fa39_3(s38[4],c38[4],andpr41[3],c39[4],s39[3]);


full_add fa39_4(s38[5],c38[5],andpr41[4],c39[5],s39[4]);


full_add fa39_5(s38[6],c38[6],andpr41[5],c39[6],s39[5]);


full_add fa39_6(s38[7],c38[7],andpr41[6],c39[7],s39[6]);


full_add fa39_7(s38[8],c38[8],andpr41[7],c39[8],s39[7]);


full_add fa39_8(s38[9],c38[9],andpr41[8],c39[9],s39[8]);


full_add fa39_9(s38[10],c38[10],andpr41[9],c39[10],s39[9]);


full_add fa39_10(s38[11],c38[11],andpr41[10],c39[11],s39[10]);


full_add fa39_11(s38[12],c38[12],andpr41[11],c39[12],s39[11]);


full_add fa39_12(s38[13],c38[13],andpr41[12],c39[13],s39[12]);


full_add fa39_13(s38[14],c38[14],andpr41[13],c39[14],s39[13]);


full_add fa39_14(s38[15],c38[15],andpr41[14],c39[15],s39[14]);


full_add fa39_15(s38[16],c38[16],andpr41[15],c39[16],s39[15]);


full_add fa39_16(s38[17],c38[17],andpr41[16],c39[17],s39[16]);


full_add fa39_17(s38[18],c38[18],andpr41[17],c39[18],s39[17]);


full_add fa39_18(s38[19],c38[19],andpr41[18],c39[19],s39[18]);


full_add fa39_19(s38[20],c38[20],andpr41[19],c39[20],s39[19]);


full_add fa39_20(s38[21],c38[21],andpr41[20],c39[21],s39[20]);


full_add fa39_21(s38[22],c38[22],andpr41[21],c39[22],s39[21]);


full_add fa39_22(s38[23],c38[23],andpr41[22],c39[23],s39[22]);


full_add fa39_23(s38[24],c38[24],andpr41[23],c39[24],s39[23]);


full_add fa39_24(s38[25],c38[25],andpr41[24],c39[25],s39[24]);


full_add fa39_25(s38[26],c38[26],andpr41[25],c39[26],s39[25]);


full_add fa39_26(s38[27],c38[27],andpr41[26],c39[27],s39[26]);


full_add fa39_27(s38[28],c38[28],andpr41[27],c39[28],s39[27]);


full_add fa39_28(s38[29],c38[29],andpr41[28],c39[29],s39[28]);


full_add fa39_29(s38[30],c38[30],andpr41[29],c39[30],s39[29]);


full_add fa39_30(s38[31],c38[31],andpr41[30],c39[31],s39[30]);


full_add fa39_31(s38[32],c38[32],andpr41[31],c39[32],s39[31]);


full_add fa39_32(s38[33],c38[33],andpr41[32],c39[33],s39[32]);


full_add fa39_33(s38[34],c38[34],andpr41[33],c39[34],s39[33]);


full_add fa39_34(s38[35],c38[35],andpr41[34],c39[35],s39[34]);


full_add fa39_35(s38[36],c38[36],andpr41[35],c39[36],s39[35]);


full_add fa39_36(s38[37],c38[37],andpr41[36],c39[37],s39[36]);


full_add fa39_37(s38[38],c38[38],andpr41[37],c39[38],s39[37]);


full_add fa39_38(s38[39],c38[39],andpr41[38],c39[39],s39[38]);


full_add fa39_39(s38[40],c38[40],andpr41[39],c39[40],s39[39]);


full_add fa39_40(s38[41],c38[41],andpr41[40],c39[41],s39[40]);


full_add fa39_41(s38[42],c38[42],andpr41[41],c39[42],s39[41]);


full_add fa39_42(s38[43],c38[43],andpr41[42],c39[43],s39[42]);


full_add fa39_43(s38[44],c38[44],andpr41[43],c39[44],s39[43]);


full_add fa39_44(s38[45],c38[45],andpr41[44],c39[45],s39[44]);


full_add fa39_45(s38[46],c38[46],andpr41[45],c39[46],s39[45]);


full_add fa39_46(s38[47],c38[47],andpr41[46],c39[47],s39[46]);


full_add fa39_47(s38[48],c38[48],andpr41[47],c39[48],s39[47]);


full_add fa39_48(s38[49],c38[49],andpr41[48],c39[49],s39[48]);


full_add fa39_49(s38[50],c38[50],andpr41[49],c39[50],s39[49]);


full_add fa39_50(s38[51],c38[51],andpr41[50],c39[51],s39[50]);


full_add fa39_51(s38[52],c38[52],andpr41[51],c39[52],s39[51]);


full_add fa39_52(s38[53],c38[53],andpr41[52],c39[53],s39[52]);


full_add fa39_53(s38[54],c38[54],andpr41[53],c39[54],s39[53]);


full_add fa39_54(s38[55],c38[55],andpr41[54],c39[55],s39[54]);


full_add fa39_55(s38[56],c38[56],andpr41[55],c39[56],s39[55]);


full_add fa39_56(s38[57],c38[57],andpr41[56],c39[57],s39[56]);


full_add fa39_57(s38[58],c38[58],andpr41[57],c39[58],s39[57]);


full_add fa39_58(s38[59],c38[59],andpr41[58],c39[59],s39[58]);


full_add fa39_59(s38[60],c38[60],andpr41[59],c39[60],s39[59]);


full_add fa39_60(s38[61],c38[61],andpr41[60],c39[61],s39[60]);


full_add fa39_61(s38[62],c38[62],andpr41[61],c39[62],s39[61]);


full_add fa39_62(si[39],c38[63],andpr41[62],c39[63],s39[62]);



half_adder ha40(s39[0],c39[0],c40[0],p[40]);


full_add fa40_0(s39[1],c39[1],andpr42[0],c40[1],s40[0]);


full_add fa40_1(s39[2],c39[2],andpr42[1],c40[2],s40[1]);


full_add fa40_2(s39[3],c39[3],andpr42[2],c40[3],s40[2]);


full_add fa40_3(s39[4],c39[4],andpr42[3],c40[4],s40[3]);


full_add fa40_4(s39[5],c39[5],andpr42[4],c40[5],s40[4]);


full_add fa40_5(s39[6],c39[6],andpr42[5],c40[6],s40[5]);


full_add fa40_6(s39[7],c39[7],andpr42[6],c40[7],s40[6]);


full_add fa40_7(s39[8],c39[8],andpr42[7],c40[8],s40[7]);


full_add fa40_8(s39[9],c39[9],andpr42[8],c40[9],s40[8]);


full_add fa40_9(s39[10],c39[10],andpr42[9],c40[10],s40[9]);


full_add fa40_10(s39[11],c39[11],andpr42[10],c40[11],s40[10]);


full_add fa40_11(s39[12],c39[12],andpr42[11],c40[12],s40[11]);


full_add fa40_12(s39[13],c39[13],andpr42[12],c40[13],s40[12]);


full_add fa40_13(s39[14],c39[14],andpr42[13],c40[14],s40[13]);


full_add fa40_14(s39[15],c39[15],andpr42[14],c40[15],s40[14]);


full_add fa40_15(s39[16],c39[16],andpr42[15],c40[16],s40[15]);


full_add fa40_16(s39[17],c39[17],andpr42[16],c40[17],s40[16]);


full_add fa40_17(s39[18],c39[18],andpr42[17],c40[18],s40[17]);


full_add fa40_18(s39[19],c39[19],andpr42[18],c40[19],s40[18]);


full_add fa40_19(s39[20],c39[20],andpr42[19],c40[20],s40[19]);


full_add fa40_20(s39[21],c39[21],andpr42[20],c40[21],s40[20]);


full_add fa40_21(s39[22],c39[22],andpr42[21],c40[22],s40[21]);


full_add fa40_22(s39[23],c39[23],andpr42[22],c40[23],s40[22]);


full_add fa40_23(s39[24],c39[24],andpr42[23],c40[24],s40[23]);


full_add fa40_24(s39[25],c39[25],andpr42[24],c40[25],s40[24]);


full_add fa40_25(s39[26],c39[26],andpr42[25],c40[26],s40[25]);


full_add fa40_26(s39[27],c39[27],andpr42[26],c40[27],s40[26]);


full_add fa40_27(s39[28],c39[28],andpr42[27],c40[28],s40[27]);


full_add fa40_28(s39[29],c39[29],andpr42[28],c40[29],s40[28]);


full_add fa40_29(s39[30],c39[30],andpr42[29],c40[30],s40[29]);


full_add fa40_30(s39[31],c39[31],andpr42[30],c40[31],s40[30]);


full_add fa40_31(s39[32],c39[32],andpr42[31],c40[32],s40[31]);


full_add fa40_32(s39[33],c39[33],andpr42[32],c40[33],s40[32]);


full_add fa40_33(s39[34],c39[34],andpr42[33],c40[34],s40[33]);


full_add fa40_34(s39[35],c39[35],andpr42[34],c40[35],s40[34]);


full_add fa40_35(s39[36],c39[36],andpr42[35],c40[36],s40[35]);


full_add fa40_36(s39[37],c39[37],andpr42[36],c40[37],s40[36]);


full_add fa40_37(s39[38],c39[38],andpr42[37],c40[38],s40[37]);


full_add fa40_38(s39[39],c39[39],andpr42[38],c40[39],s40[38]);


full_add fa40_39(s39[40],c39[40],andpr42[39],c40[40],s40[39]);


full_add fa40_40(s39[41],c39[41],andpr42[40],c40[41],s40[40]);


full_add fa40_41(s39[42],c39[42],andpr42[41],c40[42],s40[41]);


full_add fa40_42(s39[43],c39[43],andpr42[42],c40[43],s40[42]);


full_add fa40_43(s39[44],c39[44],andpr42[43],c40[44],s40[43]);


full_add fa40_44(s39[45],c39[45],andpr42[44],c40[45],s40[44]);


full_add fa40_45(s39[46],c39[46],andpr42[45],c40[46],s40[45]);


full_add fa40_46(s39[47],c39[47],andpr42[46],c40[47],s40[46]);


full_add fa40_47(s39[48],c39[48],andpr42[47],c40[48],s40[47]);


full_add fa40_48(s39[49],c39[49],andpr42[48],c40[49],s40[48]);


full_add fa40_49(s39[50],c39[50],andpr42[49],c40[50],s40[49]);


full_add fa40_50(s39[51],c39[51],andpr42[50],c40[51],s40[50]);


full_add fa40_51(s39[52],c39[52],andpr42[51],c40[52],s40[51]);


full_add fa40_52(s39[53],c39[53],andpr42[52],c40[53],s40[52]);


full_add fa40_53(s39[54],c39[54],andpr42[53],c40[54],s40[53]);


full_add fa40_54(s39[55],c39[55],andpr42[54],c40[55],s40[54]);


full_add fa40_55(s39[56],c39[56],andpr42[55],c40[56],s40[55]);


full_add fa40_56(s39[57],c39[57],andpr42[56],c40[57],s40[56]);


full_add fa40_57(s39[58],c39[58],andpr42[57],c40[58],s40[57]);


full_add fa40_58(s39[59],c39[59],andpr42[58],c40[59],s40[58]);


full_add fa40_59(s39[60],c39[60],andpr42[59],c40[60],s40[59]);


full_add fa40_60(s39[61],c39[61],andpr42[60],c40[61],s40[60]);


full_add fa40_61(s39[62],c39[62],andpr42[61],c40[62],s40[61]);


full_add fa40_62(si[40],c39[63],andpr42[62],c40[63],s40[62]);



half_adder ha41(s40[0],c40[0],c41[0],p[41]);


full_add fa41_0(s40[1],c40[1],andpr43[0],c41[1],s41[0]);


full_add fa41_1(s40[2],c40[2],andpr43[1],c41[2],s41[1]);


full_add fa41_2(s40[3],c40[3],andpr43[2],c41[3],s41[2]);


full_add fa41_3(s40[4],c40[4],andpr43[3],c41[4],s41[3]);


full_add fa41_4(s40[5],c40[5],andpr43[4],c41[5],s41[4]);


full_add fa41_5(s40[6],c40[6],andpr43[5],c41[6],s41[5]);


full_add fa41_6(s40[7],c40[7],andpr43[6],c41[7],s41[6]);


full_add fa41_7(s40[8],c40[8],andpr43[7],c41[8],s41[7]);


full_add fa41_8(s40[9],c40[9],andpr43[8],c41[9],s41[8]);


full_add fa41_9(s40[10],c40[10],andpr43[9],c41[10],s41[9]);


full_add fa41_10(s40[11],c40[11],andpr43[10],c41[11],s41[10]);


full_add fa41_11(s40[12],c40[12],andpr43[11],c41[12],s41[11]);


full_add fa41_12(s40[13],c40[13],andpr43[12],c41[13],s41[12]);


full_add fa41_13(s40[14],c40[14],andpr43[13],c41[14],s41[13]);


full_add fa41_14(s40[15],c40[15],andpr43[14],c41[15],s41[14]);


full_add fa41_15(s40[16],c40[16],andpr43[15],c41[16],s41[15]);


full_add fa41_16(s40[17],c40[17],andpr43[16],c41[17],s41[16]);


full_add fa41_17(s40[18],c40[18],andpr43[17],c41[18],s41[17]);


full_add fa41_18(s40[19],c40[19],andpr43[18],c41[19],s41[18]);


full_add fa41_19(s40[20],c40[20],andpr43[19],c41[20],s41[19]);


full_add fa41_20(s40[21],c40[21],andpr43[20],c41[21],s41[20]);


full_add fa41_21(s40[22],c40[22],andpr43[21],c41[22],s41[21]);


full_add fa41_22(s40[23],c40[23],andpr43[22],c41[23],s41[22]);


full_add fa41_23(s40[24],c40[24],andpr43[23],c41[24],s41[23]);


full_add fa41_24(s40[25],c40[25],andpr43[24],c41[25],s41[24]);


full_add fa41_25(s40[26],c40[26],andpr43[25],c41[26],s41[25]);


full_add fa41_26(s40[27],c40[27],andpr43[26],c41[27],s41[26]);


full_add fa41_27(s40[28],c40[28],andpr43[27],c41[28],s41[27]);


full_add fa41_28(s40[29],c40[29],andpr43[28],c41[29],s41[28]);


full_add fa41_29(s40[30],c40[30],andpr43[29],c41[30],s41[29]);


full_add fa41_30(s40[31],c40[31],andpr43[30],c41[31],s41[30]);


full_add fa41_31(s40[32],c40[32],andpr43[31],c41[32],s41[31]);


full_add fa41_32(s40[33],c40[33],andpr43[32],c41[33],s41[32]);


full_add fa41_33(s40[34],c40[34],andpr43[33],c41[34],s41[33]);


full_add fa41_34(s40[35],c40[35],andpr43[34],c41[35],s41[34]);


full_add fa41_35(s40[36],c40[36],andpr43[35],c41[36],s41[35]);


full_add fa41_36(s40[37],c40[37],andpr43[36],c41[37],s41[36]);


full_add fa41_37(s40[38],c40[38],andpr43[37],c41[38],s41[37]);


full_add fa41_38(s40[39],c40[39],andpr43[38],c41[39],s41[38]);


full_add fa41_39(s40[40],c40[40],andpr43[39],c41[40],s41[39]);


full_add fa41_40(s40[41],c40[41],andpr43[40],c41[41],s41[40]);


full_add fa41_41(s40[42],c40[42],andpr43[41],c41[42],s41[41]);


full_add fa41_42(s40[43],c40[43],andpr43[42],c41[43],s41[42]);


full_add fa41_43(s40[44],c40[44],andpr43[43],c41[44],s41[43]);


full_add fa41_44(s40[45],c40[45],andpr43[44],c41[45],s41[44]);


full_add fa41_45(s40[46],c40[46],andpr43[45],c41[46],s41[45]);


full_add fa41_46(s40[47],c40[47],andpr43[46],c41[47],s41[46]);


full_add fa41_47(s40[48],c40[48],andpr43[47],c41[48],s41[47]);


full_add fa41_48(s40[49],c40[49],andpr43[48],c41[49],s41[48]);


full_add fa41_49(s40[50],c40[50],andpr43[49],c41[50],s41[49]);


full_add fa41_50(s40[51],c40[51],andpr43[50],c41[51],s41[50]);


full_add fa41_51(s40[52],c40[52],andpr43[51],c41[52],s41[51]);


full_add fa41_52(s40[53],c40[53],andpr43[52],c41[53],s41[52]);


full_add fa41_53(s40[54],c40[54],andpr43[53],c41[54],s41[53]);


full_add fa41_54(s40[55],c40[55],andpr43[54],c41[55],s41[54]);


full_add fa41_55(s40[56],c40[56],andpr43[55],c41[56],s41[55]);


full_add fa41_56(s40[57],c40[57],andpr43[56],c41[57],s41[56]);


full_add fa41_57(s40[58],c40[58],andpr43[57],c41[58],s41[57]);


full_add fa41_58(s40[59],c40[59],andpr43[58],c41[59],s41[58]);


full_add fa41_59(s40[60],c40[60],andpr43[59],c41[60],s41[59]);


full_add fa41_60(s40[61],c40[61],andpr43[60],c41[61],s41[60]);


full_add fa41_61(s40[62],c40[62],andpr43[61],c41[62],s41[61]);


full_add fa41_62(si[41],c40[63],andpr43[62],c41[63],s41[62]);



half_adder ha42(s41[0],c41[0],c42[0],p[42]);


full_add fa42_0(s41[1],c41[1],andpr44[0],c42[1],s42[0]);


full_add fa42_1(s41[2],c41[2],andpr44[1],c42[2],s42[1]);


full_add fa42_2(s41[3],c41[3],andpr44[2],c42[3],s42[2]);


full_add fa42_3(s41[4],c41[4],andpr44[3],c42[4],s42[3]);


full_add fa42_4(s41[5],c41[5],andpr44[4],c42[5],s42[4]);


full_add fa42_5(s41[6],c41[6],andpr44[5],c42[6],s42[5]);


full_add fa42_6(s41[7],c41[7],andpr44[6],c42[7],s42[6]);


full_add fa42_7(s41[8],c41[8],andpr44[7],c42[8],s42[7]);


full_add fa42_8(s41[9],c41[9],andpr44[8],c42[9],s42[8]);


full_add fa42_9(s41[10],c41[10],andpr44[9],c42[10],s42[9]);


full_add fa42_10(s41[11],c41[11],andpr44[10],c42[11],s42[10]);


full_add fa42_11(s41[12],c41[12],andpr44[11],c42[12],s42[11]);


full_add fa42_12(s41[13],c41[13],andpr44[12],c42[13],s42[12]);


full_add fa42_13(s41[14],c41[14],andpr44[13],c42[14],s42[13]);


full_add fa42_14(s41[15],c41[15],andpr44[14],c42[15],s42[14]);


full_add fa42_15(s41[16],c41[16],andpr44[15],c42[16],s42[15]);


full_add fa42_16(s41[17],c41[17],andpr44[16],c42[17],s42[16]);


full_add fa42_17(s41[18],c41[18],andpr44[17],c42[18],s42[17]);


full_add fa42_18(s41[19],c41[19],andpr44[18],c42[19],s42[18]);


full_add fa42_19(s41[20],c41[20],andpr44[19],c42[20],s42[19]);


full_add fa42_20(s41[21],c41[21],andpr44[20],c42[21],s42[20]);


full_add fa42_21(s41[22],c41[22],andpr44[21],c42[22],s42[21]);


full_add fa42_22(s41[23],c41[23],andpr44[22],c42[23],s42[22]);


full_add fa42_23(s41[24],c41[24],andpr44[23],c42[24],s42[23]);


full_add fa42_24(s41[25],c41[25],andpr44[24],c42[25],s42[24]);


full_add fa42_25(s41[26],c41[26],andpr44[25],c42[26],s42[25]);


full_add fa42_26(s41[27],c41[27],andpr44[26],c42[27],s42[26]);


full_add fa42_27(s41[28],c41[28],andpr44[27],c42[28],s42[27]);


full_add fa42_28(s41[29],c41[29],andpr44[28],c42[29],s42[28]);


full_add fa42_29(s41[30],c41[30],andpr44[29],c42[30],s42[29]);


full_add fa42_30(s41[31],c41[31],andpr44[30],c42[31],s42[30]);


full_add fa42_31(s41[32],c41[32],andpr44[31],c42[32],s42[31]);


full_add fa42_32(s41[33],c41[33],andpr44[32],c42[33],s42[32]);


full_add fa42_33(s41[34],c41[34],andpr44[33],c42[34],s42[33]);


full_add fa42_34(s41[35],c41[35],andpr44[34],c42[35],s42[34]);


full_add fa42_35(s41[36],c41[36],andpr44[35],c42[36],s42[35]);


full_add fa42_36(s41[37],c41[37],andpr44[36],c42[37],s42[36]);


full_add fa42_37(s41[38],c41[38],andpr44[37],c42[38],s42[37]);


full_add fa42_38(s41[39],c41[39],andpr44[38],c42[39],s42[38]);


full_add fa42_39(s41[40],c41[40],andpr44[39],c42[40],s42[39]);


full_add fa42_40(s41[41],c41[41],andpr44[40],c42[41],s42[40]);


full_add fa42_41(s41[42],c41[42],andpr44[41],c42[42],s42[41]);


full_add fa42_42(s41[43],c41[43],andpr44[42],c42[43],s42[42]);


full_add fa42_43(s41[44],c41[44],andpr44[43],c42[44],s42[43]);


full_add fa42_44(s41[45],c41[45],andpr44[44],c42[45],s42[44]);


full_add fa42_45(s41[46],c41[46],andpr44[45],c42[46],s42[45]);


full_add fa42_46(s41[47],c41[47],andpr44[46],c42[47],s42[46]);


full_add fa42_47(s41[48],c41[48],andpr44[47],c42[48],s42[47]);


full_add fa42_48(s41[49],c41[49],andpr44[48],c42[49],s42[48]);


full_add fa42_49(s41[50],c41[50],andpr44[49],c42[50],s42[49]);


full_add fa42_50(s41[51],c41[51],andpr44[50],c42[51],s42[50]);


full_add fa42_51(s41[52],c41[52],andpr44[51],c42[52],s42[51]);


full_add fa42_52(s41[53],c41[53],andpr44[52],c42[53],s42[52]);


full_add fa42_53(s41[54],c41[54],andpr44[53],c42[54],s42[53]);


full_add fa42_54(s41[55],c41[55],andpr44[54],c42[55],s42[54]);


full_add fa42_55(s41[56],c41[56],andpr44[55],c42[56],s42[55]);


full_add fa42_56(s41[57],c41[57],andpr44[56],c42[57],s42[56]);


full_add fa42_57(s41[58],c41[58],andpr44[57],c42[58],s42[57]);


full_add fa42_58(s41[59],c41[59],andpr44[58],c42[59],s42[58]);


full_add fa42_59(s41[60],c41[60],andpr44[59],c42[60],s42[59]);


full_add fa42_60(s41[61],c41[61],andpr44[60],c42[61],s42[60]);


full_add fa42_61(s41[62],c41[62],andpr44[61],c42[62],s42[61]);


full_add fa42_62(si[42],c41[63],andpr44[62],c42[63],s42[62]);



half_adder ha43(s42[0],c42[0],c43[0],p[43]);


full_add fa43_0(s42[1],c42[1],andpr45[0],c43[1],s43[0]);


full_add fa43_1(s42[2],c42[2],andpr45[1],c43[2],s43[1]);


full_add fa43_2(s42[3],c42[3],andpr45[2],c43[3],s43[2]);


full_add fa43_3(s42[4],c42[4],andpr45[3],c43[4],s43[3]);


full_add fa43_4(s42[5],c42[5],andpr45[4],c43[5],s43[4]);


full_add fa43_5(s42[6],c42[6],andpr45[5],c43[6],s43[5]);


full_add fa43_6(s42[7],c42[7],andpr45[6],c43[7],s43[6]);


full_add fa43_7(s42[8],c42[8],andpr45[7],c43[8],s43[7]);


full_add fa43_8(s42[9],c42[9],andpr45[8],c43[9],s43[8]);


full_add fa43_9(s42[10],c42[10],andpr45[9],c43[10],s43[9]);


full_add fa43_10(s42[11],c42[11],andpr45[10],c43[11],s43[10]);


full_add fa43_11(s42[12],c42[12],andpr45[11],c43[12],s43[11]);


full_add fa43_12(s42[13],c42[13],andpr45[12],c43[13],s43[12]);


full_add fa43_13(s42[14],c42[14],andpr45[13],c43[14],s43[13]);


full_add fa43_14(s42[15],c42[15],andpr45[14],c43[15],s43[14]);


full_add fa43_15(s42[16],c42[16],andpr45[15],c43[16],s43[15]);


full_add fa43_16(s42[17],c42[17],andpr45[16],c43[17],s43[16]);


full_add fa43_17(s42[18],c42[18],andpr45[17],c43[18],s43[17]);


full_add fa43_18(s42[19],c42[19],andpr45[18],c43[19],s43[18]);


full_add fa43_19(s42[20],c42[20],andpr45[19],c43[20],s43[19]);


full_add fa43_20(s42[21],c42[21],andpr45[20],c43[21],s43[20]);


full_add fa43_21(s42[22],c42[22],andpr45[21],c43[22],s43[21]);


full_add fa43_22(s42[23],c42[23],andpr45[22],c43[23],s43[22]);


full_add fa43_23(s42[24],c42[24],andpr45[23],c43[24],s43[23]);


full_add fa43_24(s42[25],c42[25],andpr45[24],c43[25],s43[24]);


full_add fa43_25(s42[26],c42[26],andpr45[25],c43[26],s43[25]);


full_add fa43_26(s42[27],c42[27],andpr45[26],c43[27],s43[26]);


full_add fa43_27(s42[28],c42[28],andpr45[27],c43[28],s43[27]);


full_add fa43_28(s42[29],c42[29],andpr45[28],c43[29],s43[28]);


full_add fa43_29(s42[30],c42[30],andpr45[29],c43[30],s43[29]);


full_add fa43_30(s42[31],c42[31],andpr45[30],c43[31],s43[30]);


full_add fa43_31(s42[32],c42[32],andpr45[31],c43[32],s43[31]);


full_add fa43_32(s42[33],c42[33],andpr45[32],c43[33],s43[32]);


full_add fa43_33(s42[34],c42[34],andpr45[33],c43[34],s43[33]);


full_add fa43_34(s42[35],c42[35],andpr45[34],c43[35],s43[34]);


full_add fa43_35(s42[36],c42[36],andpr45[35],c43[36],s43[35]);


full_add fa43_36(s42[37],c42[37],andpr45[36],c43[37],s43[36]);


full_add fa43_37(s42[38],c42[38],andpr45[37],c43[38],s43[37]);


full_add fa43_38(s42[39],c42[39],andpr45[38],c43[39],s43[38]);


full_add fa43_39(s42[40],c42[40],andpr45[39],c43[40],s43[39]);


full_add fa43_40(s42[41],c42[41],andpr45[40],c43[41],s43[40]);


full_add fa43_41(s42[42],c42[42],andpr45[41],c43[42],s43[41]);


full_add fa43_42(s42[43],c42[43],andpr45[42],c43[43],s43[42]);


full_add fa43_43(s42[44],c42[44],andpr45[43],c43[44],s43[43]);


full_add fa43_44(s42[45],c42[45],andpr45[44],c43[45],s43[44]);


full_add fa43_45(s42[46],c42[46],andpr45[45],c43[46],s43[45]);


full_add fa43_46(s42[47],c42[47],andpr45[46],c43[47],s43[46]);


full_add fa43_47(s42[48],c42[48],andpr45[47],c43[48],s43[47]);


full_add fa43_48(s42[49],c42[49],andpr45[48],c43[49],s43[48]);


full_add fa43_49(s42[50],c42[50],andpr45[49],c43[50],s43[49]);


full_add fa43_50(s42[51],c42[51],andpr45[50],c43[51],s43[50]);


full_add fa43_51(s42[52],c42[52],andpr45[51],c43[52],s43[51]);


full_add fa43_52(s42[53],c42[53],andpr45[52],c43[53],s43[52]);


full_add fa43_53(s42[54],c42[54],andpr45[53],c43[54],s43[53]);


full_add fa43_54(s42[55],c42[55],andpr45[54],c43[55],s43[54]);


full_add fa43_55(s42[56],c42[56],andpr45[55],c43[56],s43[55]);


full_add fa43_56(s42[57],c42[57],andpr45[56],c43[57],s43[56]);


full_add fa43_57(s42[58],c42[58],andpr45[57],c43[58],s43[57]);


full_add fa43_58(s42[59],c42[59],andpr45[58],c43[59],s43[58]);


full_add fa43_59(s42[60],c42[60],andpr45[59],c43[60],s43[59]);


full_add fa43_60(s42[61],c42[61],andpr45[60],c43[61],s43[60]);


full_add fa43_61(s42[62],c42[62],andpr45[61],c43[62],s43[61]);


full_add fa43_62(si[43],c42[63],andpr45[62],c43[63],s43[62]);



half_adder ha44(s43[0],c43[0],c44[0],p[44]);


full_add fa44_0(s43[1],c43[1],andpr46[0],c44[1],s44[0]);


full_add fa44_1(s43[2],c43[2],andpr46[1],c44[2],s44[1]);


full_add fa44_2(s43[3],c43[3],andpr46[2],c44[3],s44[2]);


full_add fa44_3(s43[4],c43[4],andpr46[3],c44[4],s44[3]);


full_add fa44_4(s43[5],c43[5],andpr46[4],c44[5],s44[4]);


full_add fa44_5(s43[6],c43[6],andpr46[5],c44[6],s44[5]);


full_add fa44_6(s43[7],c43[7],andpr46[6],c44[7],s44[6]);


full_add fa44_7(s43[8],c43[8],andpr46[7],c44[8],s44[7]);


full_add fa44_8(s43[9],c43[9],andpr46[8],c44[9],s44[8]);


full_add fa44_9(s43[10],c43[10],andpr46[9],c44[10],s44[9]);


full_add fa44_10(s43[11],c43[11],andpr46[10],c44[11],s44[10]);


full_add fa44_11(s43[12],c43[12],andpr46[11],c44[12],s44[11]);


full_add fa44_12(s43[13],c43[13],andpr46[12],c44[13],s44[12]);


full_add fa44_13(s43[14],c43[14],andpr46[13],c44[14],s44[13]);


full_add fa44_14(s43[15],c43[15],andpr46[14],c44[15],s44[14]);


full_add fa44_15(s43[16],c43[16],andpr46[15],c44[16],s44[15]);


full_add fa44_16(s43[17],c43[17],andpr46[16],c44[17],s44[16]);


full_add fa44_17(s43[18],c43[18],andpr46[17],c44[18],s44[17]);


full_add fa44_18(s43[19],c43[19],andpr46[18],c44[19],s44[18]);


full_add fa44_19(s43[20],c43[20],andpr46[19],c44[20],s44[19]);


full_add fa44_20(s43[21],c43[21],andpr46[20],c44[21],s44[20]);


full_add fa44_21(s43[22],c43[22],andpr46[21],c44[22],s44[21]);


full_add fa44_22(s43[23],c43[23],andpr46[22],c44[23],s44[22]);


full_add fa44_23(s43[24],c43[24],andpr46[23],c44[24],s44[23]);


full_add fa44_24(s43[25],c43[25],andpr46[24],c44[25],s44[24]);


full_add fa44_25(s43[26],c43[26],andpr46[25],c44[26],s44[25]);


full_add fa44_26(s43[27],c43[27],andpr46[26],c44[27],s44[26]);


full_add fa44_27(s43[28],c43[28],andpr46[27],c44[28],s44[27]);


full_add fa44_28(s43[29],c43[29],andpr46[28],c44[29],s44[28]);


full_add fa44_29(s43[30],c43[30],andpr46[29],c44[30],s44[29]);


full_add fa44_30(s43[31],c43[31],andpr46[30],c44[31],s44[30]);


full_add fa44_31(s43[32],c43[32],andpr46[31],c44[32],s44[31]);


full_add fa44_32(s43[33],c43[33],andpr46[32],c44[33],s44[32]);


full_add fa44_33(s43[34],c43[34],andpr46[33],c44[34],s44[33]);


full_add fa44_34(s43[35],c43[35],andpr46[34],c44[35],s44[34]);


full_add fa44_35(s43[36],c43[36],andpr46[35],c44[36],s44[35]);


full_add fa44_36(s43[37],c43[37],andpr46[36],c44[37],s44[36]);


full_add fa44_37(s43[38],c43[38],andpr46[37],c44[38],s44[37]);


full_add fa44_38(s43[39],c43[39],andpr46[38],c44[39],s44[38]);


full_add fa44_39(s43[40],c43[40],andpr46[39],c44[40],s44[39]);


full_add fa44_40(s43[41],c43[41],andpr46[40],c44[41],s44[40]);


full_add fa44_41(s43[42],c43[42],andpr46[41],c44[42],s44[41]);


full_add fa44_42(s43[43],c43[43],andpr46[42],c44[43],s44[42]);


full_add fa44_43(s43[44],c43[44],andpr46[43],c44[44],s44[43]);


full_add fa44_44(s43[45],c43[45],andpr46[44],c44[45],s44[44]);


full_add fa44_45(s43[46],c43[46],andpr46[45],c44[46],s44[45]);


full_add fa44_46(s43[47],c43[47],andpr46[46],c44[47],s44[46]);


full_add fa44_47(s43[48],c43[48],andpr46[47],c44[48],s44[47]);


full_add fa44_48(s43[49],c43[49],andpr46[48],c44[49],s44[48]);


full_add fa44_49(s43[50],c43[50],andpr46[49],c44[50],s44[49]);


full_add fa44_50(s43[51],c43[51],andpr46[50],c44[51],s44[50]);


full_add fa44_51(s43[52],c43[52],andpr46[51],c44[52],s44[51]);


full_add fa44_52(s43[53],c43[53],andpr46[52],c44[53],s44[52]);


full_add fa44_53(s43[54],c43[54],andpr46[53],c44[54],s44[53]);


full_add fa44_54(s43[55],c43[55],andpr46[54],c44[55],s44[54]);


full_add fa44_55(s43[56],c43[56],andpr46[55],c44[56],s44[55]);


full_add fa44_56(s43[57],c43[57],andpr46[56],c44[57],s44[56]);


full_add fa44_57(s43[58],c43[58],andpr46[57],c44[58],s44[57]);


full_add fa44_58(s43[59],c43[59],andpr46[58],c44[59],s44[58]);


full_add fa44_59(s43[60],c43[60],andpr46[59],c44[60],s44[59]);


full_add fa44_60(s43[61],c43[61],andpr46[60],c44[61],s44[60]);


full_add fa44_61(s43[62],c43[62],andpr46[61],c44[62],s44[61]);


full_add fa44_62(si[44],c43[63],andpr46[62],c44[63],s44[62]);



half_adder ha45(s44[0],c44[0],c45[0],p[45]);


full_add fa45_0(s44[1],c44[1],andpr47[0],c45[1],s45[0]);


full_add fa45_1(s44[2],c44[2],andpr47[1],c45[2],s45[1]);


full_add fa45_2(s44[3],c44[3],andpr47[2],c45[3],s45[2]);


full_add fa45_3(s44[4],c44[4],andpr47[3],c45[4],s45[3]);


full_add fa45_4(s44[5],c44[5],andpr47[4],c45[5],s45[4]);


full_add fa45_5(s44[6],c44[6],andpr47[5],c45[6],s45[5]);


full_add fa45_6(s44[7],c44[7],andpr47[6],c45[7],s45[6]);


full_add fa45_7(s44[8],c44[8],andpr47[7],c45[8],s45[7]);


full_add fa45_8(s44[9],c44[9],andpr47[8],c45[9],s45[8]);


full_add fa45_9(s44[10],c44[10],andpr47[9],c45[10],s45[9]);


full_add fa45_10(s44[11],c44[11],andpr47[10],c45[11],s45[10]);


full_add fa45_11(s44[12],c44[12],andpr47[11],c45[12],s45[11]);


full_add fa45_12(s44[13],c44[13],andpr47[12],c45[13],s45[12]);


full_add fa45_13(s44[14],c44[14],andpr47[13],c45[14],s45[13]);


full_add fa45_14(s44[15],c44[15],andpr47[14],c45[15],s45[14]);


full_add fa45_15(s44[16],c44[16],andpr47[15],c45[16],s45[15]);


full_add fa45_16(s44[17],c44[17],andpr47[16],c45[17],s45[16]);


full_add fa45_17(s44[18],c44[18],andpr47[17],c45[18],s45[17]);


full_add fa45_18(s44[19],c44[19],andpr47[18],c45[19],s45[18]);


full_add fa45_19(s44[20],c44[20],andpr47[19],c45[20],s45[19]);


full_add fa45_20(s44[21],c44[21],andpr47[20],c45[21],s45[20]);


full_add fa45_21(s44[22],c44[22],andpr47[21],c45[22],s45[21]);


full_add fa45_22(s44[23],c44[23],andpr47[22],c45[23],s45[22]);


full_add fa45_23(s44[24],c44[24],andpr47[23],c45[24],s45[23]);


full_add fa45_24(s44[25],c44[25],andpr47[24],c45[25],s45[24]);


full_add fa45_25(s44[26],c44[26],andpr47[25],c45[26],s45[25]);


full_add fa45_26(s44[27],c44[27],andpr47[26],c45[27],s45[26]);


full_add fa45_27(s44[28],c44[28],andpr47[27],c45[28],s45[27]);


full_add fa45_28(s44[29],c44[29],andpr47[28],c45[29],s45[28]);


full_add fa45_29(s44[30],c44[30],andpr47[29],c45[30],s45[29]);


full_add fa45_30(s44[31],c44[31],andpr47[30],c45[31],s45[30]);


full_add fa45_31(s44[32],c44[32],andpr47[31],c45[32],s45[31]);


full_add fa45_32(s44[33],c44[33],andpr47[32],c45[33],s45[32]);


full_add fa45_33(s44[34],c44[34],andpr47[33],c45[34],s45[33]);


full_add fa45_34(s44[35],c44[35],andpr47[34],c45[35],s45[34]);


full_add fa45_35(s44[36],c44[36],andpr47[35],c45[36],s45[35]);


full_add fa45_36(s44[37],c44[37],andpr47[36],c45[37],s45[36]);


full_add fa45_37(s44[38],c44[38],andpr47[37],c45[38],s45[37]);


full_add fa45_38(s44[39],c44[39],andpr47[38],c45[39],s45[38]);


full_add fa45_39(s44[40],c44[40],andpr47[39],c45[40],s45[39]);


full_add fa45_40(s44[41],c44[41],andpr47[40],c45[41],s45[40]);


full_add fa45_41(s44[42],c44[42],andpr47[41],c45[42],s45[41]);


full_add fa45_42(s44[43],c44[43],andpr47[42],c45[43],s45[42]);


full_add fa45_43(s44[44],c44[44],andpr47[43],c45[44],s45[43]);


full_add fa45_44(s44[45],c44[45],andpr47[44],c45[45],s45[44]);


full_add fa45_45(s44[46],c44[46],andpr47[45],c45[46],s45[45]);


full_add fa45_46(s44[47],c44[47],andpr47[46],c45[47],s45[46]);


full_add fa45_47(s44[48],c44[48],andpr47[47],c45[48],s45[47]);


full_add fa45_48(s44[49],c44[49],andpr47[48],c45[49],s45[48]);


full_add fa45_49(s44[50],c44[50],andpr47[49],c45[50],s45[49]);


full_add fa45_50(s44[51],c44[51],andpr47[50],c45[51],s45[50]);


full_add fa45_51(s44[52],c44[52],andpr47[51],c45[52],s45[51]);


full_add fa45_52(s44[53],c44[53],andpr47[52],c45[53],s45[52]);


full_add fa45_53(s44[54],c44[54],andpr47[53],c45[54],s45[53]);


full_add fa45_54(s44[55],c44[55],andpr47[54],c45[55],s45[54]);


full_add fa45_55(s44[56],c44[56],andpr47[55],c45[56],s45[55]);


full_add fa45_56(s44[57],c44[57],andpr47[56],c45[57],s45[56]);


full_add fa45_57(s44[58],c44[58],andpr47[57],c45[58],s45[57]);


full_add fa45_58(s44[59],c44[59],andpr47[58],c45[59],s45[58]);


full_add fa45_59(s44[60],c44[60],andpr47[59],c45[60],s45[59]);


full_add fa45_60(s44[61],c44[61],andpr47[60],c45[61],s45[60]);


full_add fa45_61(s44[62],c44[62],andpr47[61],c45[62],s45[61]);


full_add fa45_62(si[45],c44[63],andpr47[62],c45[63],s45[62]);



half_adder ha46(s45[0],c45[0],c46[0],p[46]);


full_add fa46_0(s45[1],c45[1],andpr48[0],c46[1],s46[0]);


full_add fa46_1(s45[2],c45[2],andpr48[1],c46[2],s46[1]);


full_add fa46_2(s45[3],c45[3],andpr48[2],c46[3],s46[2]);


full_add fa46_3(s45[4],c45[4],andpr48[3],c46[4],s46[3]);


full_add fa46_4(s45[5],c45[5],andpr48[4],c46[5],s46[4]);


full_add fa46_5(s45[6],c45[6],andpr48[5],c46[6],s46[5]);


full_add fa46_6(s45[7],c45[7],andpr48[6],c46[7],s46[6]);


full_add fa46_7(s45[8],c45[8],andpr48[7],c46[8],s46[7]);


full_add fa46_8(s45[9],c45[9],andpr48[8],c46[9],s46[8]);


full_add fa46_9(s45[10],c45[10],andpr48[9],c46[10],s46[9]);


full_add fa46_10(s45[11],c45[11],andpr48[10],c46[11],s46[10]);


full_add fa46_11(s45[12],c45[12],andpr48[11],c46[12],s46[11]);


full_add fa46_12(s45[13],c45[13],andpr48[12],c46[13],s46[12]);


full_add fa46_13(s45[14],c45[14],andpr48[13],c46[14],s46[13]);


full_add fa46_14(s45[15],c45[15],andpr48[14],c46[15],s46[14]);


full_add fa46_15(s45[16],c45[16],andpr48[15],c46[16],s46[15]);


full_add fa46_16(s45[17],c45[17],andpr48[16],c46[17],s46[16]);


full_add fa46_17(s45[18],c45[18],andpr48[17],c46[18],s46[17]);


full_add fa46_18(s45[19],c45[19],andpr48[18],c46[19],s46[18]);


full_add fa46_19(s45[20],c45[20],andpr48[19],c46[20],s46[19]);


full_add fa46_20(s45[21],c45[21],andpr48[20],c46[21],s46[20]);


full_add fa46_21(s45[22],c45[22],andpr48[21],c46[22],s46[21]);


full_add fa46_22(s45[23],c45[23],andpr48[22],c46[23],s46[22]);


full_add fa46_23(s45[24],c45[24],andpr48[23],c46[24],s46[23]);


full_add fa46_24(s45[25],c45[25],andpr48[24],c46[25],s46[24]);


full_add fa46_25(s45[26],c45[26],andpr48[25],c46[26],s46[25]);


full_add fa46_26(s45[27],c45[27],andpr48[26],c46[27],s46[26]);


full_add fa46_27(s45[28],c45[28],andpr48[27],c46[28],s46[27]);


full_add fa46_28(s45[29],c45[29],andpr48[28],c46[29],s46[28]);


full_add fa46_29(s45[30],c45[30],andpr48[29],c46[30],s46[29]);


full_add fa46_30(s45[31],c45[31],andpr48[30],c46[31],s46[30]);


full_add fa46_31(s45[32],c45[32],andpr48[31],c46[32],s46[31]);


full_add fa46_32(s45[33],c45[33],andpr48[32],c46[33],s46[32]);


full_add fa46_33(s45[34],c45[34],andpr48[33],c46[34],s46[33]);


full_add fa46_34(s45[35],c45[35],andpr48[34],c46[35],s46[34]);


full_add fa46_35(s45[36],c45[36],andpr48[35],c46[36],s46[35]);


full_add fa46_36(s45[37],c45[37],andpr48[36],c46[37],s46[36]);


full_add fa46_37(s45[38],c45[38],andpr48[37],c46[38],s46[37]);


full_add fa46_38(s45[39],c45[39],andpr48[38],c46[39],s46[38]);


full_add fa46_39(s45[40],c45[40],andpr48[39],c46[40],s46[39]);


full_add fa46_40(s45[41],c45[41],andpr48[40],c46[41],s46[40]);


full_add fa46_41(s45[42],c45[42],andpr48[41],c46[42],s46[41]);


full_add fa46_42(s45[43],c45[43],andpr48[42],c46[43],s46[42]);


full_add fa46_43(s45[44],c45[44],andpr48[43],c46[44],s46[43]);


full_add fa46_44(s45[45],c45[45],andpr48[44],c46[45],s46[44]);


full_add fa46_45(s45[46],c45[46],andpr48[45],c46[46],s46[45]);


full_add fa46_46(s45[47],c45[47],andpr48[46],c46[47],s46[46]);


full_add fa46_47(s45[48],c45[48],andpr48[47],c46[48],s46[47]);


full_add fa46_48(s45[49],c45[49],andpr48[48],c46[49],s46[48]);


full_add fa46_49(s45[50],c45[50],andpr48[49],c46[50],s46[49]);


full_add fa46_50(s45[51],c45[51],andpr48[50],c46[51],s46[50]);


full_add fa46_51(s45[52],c45[52],andpr48[51],c46[52],s46[51]);


full_add fa46_52(s45[53],c45[53],andpr48[52],c46[53],s46[52]);


full_add fa46_53(s45[54],c45[54],andpr48[53],c46[54],s46[53]);


full_add fa46_54(s45[55],c45[55],andpr48[54],c46[55],s46[54]);


full_add fa46_55(s45[56],c45[56],andpr48[55],c46[56],s46[55]);


full_add fa46_56(s45[57],c45[57],andpr48[56],c46[57],s46[56]);


full_add fa46_57(s45[58],c45[58],andpr48[57],c46[58],s46[57]);


full_add fa46_58(s45[59],c45[59],andpr48[58],c46[59],s46[58]);


full_add fa46_59(s45[60],c45[60],andpr48[59],c46[60],s46[59]);


full_add fa46_60(s45[61],c45[61],andpr48[60],c46[61],s46[60]);


full_add fa46_61(s45[62],c45[62],andpr48[61],c46[62],s46[61]);


full_add fa46_62(si[46],c45[63],andpr48[62],c46[63],s46[62]);



half_adder ha47(s46[0],c46[0],c47[0],p[47]);


full_add fa47_0(s46[1],c46[1],andpr49[0],c47[1],s47[0]);


full_add fa47_1(s46[2],c46[2],andpr49[1],c47[2],s47[1]);


full_add fa47_2(s46[3],c46[3],andpr49[2],c47[3],s47[2]);


full_add fa47_3(s46[4],c46[4],andpr49[3],c47[4],s47[3]);


full_add fa47_4(s46[5],c46[5],andpr49[4],c47[5],s47[4]);


full_add fa47_5(s46[6],c46[6],andpr49[5],c47[6],s47[5]);


full_add fa47_6(s46[7],c46[7],andpr49[6],c47[7],s47[6]);


full_add fa47_7(s46[8],c46[8],andpr49[7],c47[8],s47[7]);


full_add fa47_8(s46[9],c46[9],andpr49[8],c47[9],s47[8]);


full_add fa47_9(s46[10],c46[10],andpr49[9],c47[10],s47[9]);


full_add fa47_10(s46[11],c46[11],andpr49[10],c47[11],s47[10]);


full_add fa47_11(s46[12],c46[12],andpr49[11],c47[12],s47[11]);


full_add fa47_12(s46[13],c46[13],andpr49[12],c47[13],s47[12]);


full_add fa47_13(s46[14],c46[14],andpr49[13],c47[14],s47[13]);


full_add fa47_14(s46[15],c46[15],andpr49[14],c47[15],s47[14]);


full_add fa47_15(s46[16],c46[16],andpr49[15],c47[16],s47[15]);


full_add fa47_16(s46[17],c46[17],andpr49[16],c47[17],s47[16]);


full_add fa47_17(s46[18],c46[18],andpr49[17],c47[18],s47[17]);


full_add fa47_18(s46[19],c46[19],andpr49[18],c47[19],s47[18]);


full_add fa47_19(s46[20],c46[20],andpr49[19],c47[20],s47[19]);


full_add fa47_20(s46[21],c46[21],andpr49[20],c47[21],s47[20]);


full_add fa47_21(s46[22],c46[22],andpr49[21],c47[22],s47[21]);


full_add fa47_22(s46[23],c46[23],andpr49[22],c47[23],s47[22]);


full_add fa47_23(s46[24],c46[24],andpr49[23],c47[24],s47[23]);


full_add fa47_24(s46[25],c46[25],andpr49[24],c47[25],s47[24]);


full_add fa47_25(s46[26],c46[26],andpr49[25],c47[26],s47[25]);


full_add fa47_26(s46[27],c46[27],andpr49[26],c47[27],s47[26]);


full_add fa47_27(s46[28],c46[28],andpr49[27],c47[28],s47[27]);


full_add fa47_28(s46[29],c46[29],andpr49[28],c47[29],s47[28]);


full_add fa47_29(s46[30],c46[30],andpr49[29],c47[30],s47[29]);


full_add fa47_30(s46[31],c46[31],andpr49[30],c47[31],s47[30]);


full_add fa47_31(s46[32],c46[32],andpr49[31],c47[32],s47[31]);


full_add fa47_32(s46[33],c46[33],andpr49[32],c47[33],s47[32]);


full_add fa47_33(s46[34],c46[34],andpr49[33],c47[34],s47[33]);


full_add fa47_34(s46[35],c46[35],andpr49[34],c47[35],s47[34]);


full_add fa47_35(s46[36],c46[36],andpr49[35],c47[36],s47[35]);


full_add fa47_36(s46[37],c46[37],andpr49[36],c47[37],s47[36]);


full_add fa47_37(s46[38],c46[38],andpr49[37],c47[38],s47[37]);


full_add fa47_38(s46[39],c46[39],andpr49[38],c47[39],s47[38]);


full_add fa47_39(s46[40],c46[40],andpr49[39],c47[40],s47[39]);


full_add fa47_40(s46[41],c46[41],andpr49[40],c47[41],s47[40]);


full_add fa47_41(s46[42],c46[42],andpr49[41],c47[42],s47[41]);


full_add fa47_42(s46[43],c46[43],andpr49[42],c47[43],s47[42]);


full_add fa47_43(s46[44],c46[44],andpr49[43],c47[44],s47[43]);


full_add fa47_44(s46[45],c46[45],andpr49[44],c47[45],s47[44]);


full_add fa47_45(s46[46],c46[46],andpr49[45],c47[46],s47[45]);


full_add fa47_46(s46[47],c46[47],andpr49[46],c47[47],s47[46]);


full_add fa47_47(s46[48],c46[48],andpr49[47],c47[48],s47[47]);


full_add fa47_48(s46[49],c46[49],andpr49[48],c47[49],s47[48]);


full_add fa47_49(s46[50],c46[50],andpr49[49],c47[50],s47[49]);


full_add fa47_50(s46[51],c46[51],andpr49[50],c47[51],s47[50]);


full_add fa47_51(s46[52],c46[52],andpr49[51],c47[52],s47[51]);


full_add fa47_52(s46[53],c46[53],andpr49[52],c47[53],s47[52]);


full_add fa47_53(s46[54],c46[54],andpr49[53],c47[54],s47[53]);


full_add fa47_54(s46[55],c46[55],andpr49[54],c47[55],s47[54]);


full_add fa47_55(s46[56],c46[56],andpr49[55],c47[56],s47[55]);


full_add fa47_56(s46[57],c46[57],andpr49[56],c47[57],s47[56]);


full_add fa47_57(s46[58],c46[58],andpr49[57],c47[58],s47[57]);


full_add fa47_58(s46[59],c46[59],andpr49[58],c47[59],s47[58]);


full_add fa47_59(s46[60],c46[60],andpr49[59],c47[60],s47[59]);


full_add fa47_60(s46[61],c46[61],andpr49[60],c47[61],s47[60]);


full_add fa47_61(s46[62],c46[62],andpr49[61],c47[62],s47[61]);


full_add fa47_62(si[47],c46[63],andpr49[62],c47[63],s47[62]);



half_adder ha48(s47[0],c47[0],c48[0],p[48]);


full_add fa48_0(s47[1],c47[1],andpr50[0],c48[1],s48[0]);


full_add fa48_1(s47[2],c47[2],andpr50[1],c48[2],s48[1]);


full_add fa48_2(s47[3],c47[3],andpr50[2],c48[3],s48[2]);


full_add fa48_3(s47[4],c47[4],andpr50[3],c48[4],s48[3]);


full_add fa48_4(s47[5],c47[5],andpr50[4],c48[5],s48[4]);


full_add fa48_5(s47[6],c47[6],andpr50[5],c48[6],s48[5]);


full_add fa48_6(s47[7],c47[7],andpr50[6],c48[7],s48[6]);


full_add fa48_7(s47[8],c47[8],andpr50[7],c48[8],s48[7]);


full_add fa48_8(s47[9],c47[9],andpr50[8],c48[9],s48[8]);


full_add fa48_9(s47[10],c47[10],andpr50[9],c48[10],s48[9]);


full_add fa48_10(s47[11],c47[11],andpr50[10],c48[11],s48[10]);


full_add fa48_11(s47[12],c47[12],andpr50[11],c48[12],s48[11]);


full_add fa48_12(s47[13],c47[13],andpr50[12],c48[13],s48[12]);


full_add fa48_13(s47[14],c47[14],andpr50[13],c48[14],s48[13]);


full_add fa48_14(s47[15],c47[15],andpr50[14],c48[15],s48[14]);


full_add fa48_15(s47[16],c47[16],andpr50[15],c48[16],s48[15]);


full_add fa48_16(s47[17],c47[17],andpr50[16],c48[17],s48[16]);


full_add fa48_17(s47[18],c47[18],andpr50[17],c48[18],s48[17]);


full_add fa48_18(s47[19],c47[19],andpr50[18],c48[19],s48[18]);


full_add fa48_19(s47[20],c47[20],andpr50[19],c48[20],s48[19]);


full_add fa48_20(s47[21],c47[21],andpr50[20],c48[21],s48[20]);


full_add fa48_21(s47[22],c47[22],andpr50[21],c48[22],s48[21]);


full_add fa48_22(s47[23],c47[23],andpr50[22],c48[23],s48[22]);


full_add fa48_23(s47[24],c47[24],andpr50[23],c48[24],s48[23]);


full_add fa48_24(s47[25],c47[25],andpr50[24],c48[25],s48[24]);


full_add fa48_25(s47[26],c47[26],andpr50[25],c48[26],s48[25]);


full_add fa48_26(s47[27],c47[27],andpr50[26],c48[27],s48[26]);


full_add fa48_27(s47[28],c47[28],andpr50[27],c48[28],s48[27]);


full_add fa48_28(s47[29],c47[29],andpr50[28],c48[29],s48[28]);


full_add fa48_29(s47[30],c47[30],andpr50[29],c48[30],s48[29]);


full_add fa48_30(s47[31],c47[31],andpr50[30],c48[31],s48[30]);


full_add fa48_31(s47[32],c47[32],andpr50[31],c48[32],s48[31]);


full_add fa48_32(s47[33],c47[33],andpr50[32],c48[33],s48[32]);


full_add fa48_33(s47[34],c47[34],andpr50[33],c48[34],s48[33]);


full_add fa48_34(s47[35],c47[35],andpr50[34],c48[35],s48[34]);


full_add fa48_35(s47[36],c47[36],andpr50[35],c48[36],s48[35]);


full_add fa48_36(s47[37],c47[37],andpr50[36],c48[37],s48[36]);


full_add fa48_37(s47[38],c47[38],andpr50[37],c48[38],s48[37]);


full_add fa48_38(s47[39],c47[39],andpr50[38],c48[39],s48[38]);


full_add fa48_39(s47[40],c47[40],andpr50[39],c48[40],s48[39]);


full_add fa48_40(s47[41],c47[41],andpr50[40],c48[41],s48[40]);


full_add fa48_41(s47[42],c47[42],andpr50[41],c48[42],s48[41]);


full_add fa48_42(s47[43],c47[43],andpr50[42],c48[43],s48[42]);


full_add fa48_43(s47[44],c47[44],andpr50[43],c48[44],s48[43]);


full_add fa48_44(s47[45],c47[45],andpr50[44],c48[45],s48[44]);


full_add fa48_45(s47[46],c47[46],andpr50[45],c48[46],s48[45]);


full_add fa48_46(s47[47],c47[47],andpr50[46],c48[47],s48[46]);


full_add fa48_47(s47[48],c47[48],andpr50[47],c48[48],s48[47]);


full_add fa48_48(s47[49],c47[49],andpr50[48],c48[49],s48[48]);


full_add fa48_49(s47[50],c47[50],andpr50[49],c48[50],s48[49]);


full_add fa48_50(s47[51],c47[51],andpr50[50],c48[51],s48[50]);


full_add fa48_51(s47[52],c47[52],andpr50[51],c48[52],s48[51]);


full_add fa48_52(s47[53],c47[53],andpr50[52],c48[53],s48[52]);


full_add fa48_53(s47[54],c47[54],andpr50[53],c48[54],s48[53]);


full_add fa48_54(s47[55],c47[55],andpr50[54],c48[55],s48[54]);


full_add fa48_55(s47[56],c47[56],andpr50[55],c48[56],s48[55]);


full_add fa48_56(s47[57],c47[57],andpr50[56],c48[57],s48[56]);


full_add fa48_57(s47[58],c47[58],andpr50[57],c48[58],s48[57]);


full_add fa48_58(s47[59],c47[59],andpr50[58],c48[59],s48[58]);


full_add fa48_59(s47[60],c47[60],andpr50[59],c48[60],s48[59]);


full_add fa48_60(s47[61],c47[61],andpr50[60],c48[61],s48[60]);


full_add fa48_61(s47[62],c47[62],andpr50[61],c48[62],s48[61]);


full_add fa48_62(si[48],c47[63],andpr50[62],c48[63],s48[62]);



half_adder ha49(s48[0],c48[0],c49[0],p[49]);


full_add fa49_0(s48[1],c48[1],andpr51[0],c49[1],s49[0]);


full_add fa49_1(s48[2],c48[2],andpr51[1],c49[2],s49[1]);


full_add fa49_2(s48[3],c48[3],andpr51[2],c49[3],s49[2]);


full_add fa49_3(s48[4],c48[4],andpr51[3],c49[4],s49[3]);


full_add fa49_4(s48[5],c48[5],andpr51[4],c49[5],s49[4]);


full_add fa49_5(s48[6],c48[6],andpr51[5],c49[6],s49[5]);


full_add fa49_6(s48[7],c48[7],andpr51[6],c49[7],s49[6]);


full_add fa49_7(s48[8],c48[8],andpr51[7],c49[8],s49[7]);


full_add fa49_8(s48[9],c48[9],andpr51[8],c49[9],s49[8]);


full_add fa49_9(s48[10],c48[10],andpr51[9],c49[10],s49[9]);


full_add fa49_10(s48[11],c48[11],andpr51[10],c49[11],s49[10]);


full_add fa49_11(s48[12],c48[12],andpr51[11],c49[12],s49[11]);


full_add fa49_12(s48[13],c48[13],andpr51[12],c49[13],s49[12]);


full_add fa49_13(s48[14],c48[14],andpr51[13],c49[14],s49[13]);


full_add fa49_14(s48[15],c48[15],andpr51[14],c49[15],s49[14]);


full_add fa49_15(s48[16],c48[16],andpr51[15],c49[16],s49[15]);


full_add fa49_16(s48[17],c48[17],andpr51[16],c49[17],s49[16]);


full_add fa49_17(s48[18],c48[18],andpr51[17],c49[18],s49[17]);


full_add fa49_18(s48[19],c48[19],andpr51[18],c49[19],s49[18]);


full_add fa49_19(s48[20],c48[20],andpr51[19],c49[20],s49[19]);


full_add fa49_20(s48[21],c48[21],andpr51[20],c49[21],s49[20]);


full_add fa49_21(s48[22],c48[22],andpr51[21],c49[22],s49[21]);


full_add fa49_22(s48[23],c48[23],andpr51[22],c49[23],s49[22]);


full_add fa49_23(s48[24],c48[24],andpr51[23],c49[24],s49[23]);


full_add fa49_24(s48[25],c48[25],andpr51[24],c49[25],s49[24]);


full_add fa49_25(s48[26],c48[26],andpr51[25],c49[26],s49[25]);


full_add fa49_26(s48[27],c48[27],andpr51[26],c49[27],s49[26]);


full_add fa49_27(s48[28],c48[28],andpr51[27],c49[28],s49[27]);


full_add fa49_28(s48[29],c48[29],andpr51[28],c49[29],s49[28]);


full_add fa49_29(s48[30],c48[30],andpr51[29],c49[30],s49[29]);


full_add fa49_30(s48[31],c48[31],andpr51[30],c49[31],s49[30]);


full_add fa49_31(s48[32],c48[32],andpr51[31],c49[32],s49[31]);


full_add fa49_32(s48[33],c48[33],andpr51[32],c49[33],s49[32]);


full_add fa49_33(s48[34],c48[34],andpr51[33],c49[34],s49[33]);


full_add fa49_34(s48[35],c48[35],andpr51[34],c49[35],s49[34]);


full_add fa49_35(s48[36],c48[36],andpr51[35],c49[36],s49[35]);


full_add fa49_36(s48[37],c48[37],andpr51[36],c49[37],s49[36]);


full_add fa49_37(s48[38],c48[38],andpr51[37],c49[38],s49[37]);


full_add fa49_38(s48[39],c48[39],andpr51[38],c49[39],s49[38]);


full_add fa49_39(s48[40],c48[40],andpr51[39],c49[40],s49[39]);


full_add fa49_40(s48[41],c48[41],andpr51[40],c49[41],s49[40]);


full_add fa49_41(s48[42],c48[42],andpr51[41],c49[42],s49[41]);


full_add fa49_42(s48[43],c48[43],andpr51[42],c49[43],s49[42]);


full_add fa49_43(s48[44],c48[44],andpr51[43],c49[44],s49[43]);


full_add fa49_44(s48[45],c48[45],andpr51[44],c49[45],s49[44]);


full_add fa49_45(s48[46],c48[46],andpr51[45],c49[46],s49[45]);


full_add fa49_46(s48[47],c48[47],andpr51[46],c49[47],s49[46]);


full_add fa49_47(s48[48],c48[48],andpr51[47],c49[48],s49[47]);


full_add fa49_48(s48[49],c48[49],andpr51[48],c49[49],s49[48]);


full_add fa49_49(s48[50],c48[50],andpr51[49],c49[50],s49[49]);


full_add fa49_50(s48[51],c48[51],andpr51[50],c49[51],s49[50]);


full_add fa49_51(s48[52],c48[52],andpr51[51],c49[52],s49[51]);


full_add fa49_52(s48[53],c48[53],andpr51[52],c49[53],s49[52]);


full_add fa49_53(s48[54],c48[54],andpr51[53],c49[54],s49[53]);


full_add fa49_54(s48[55],c48[55],andpr51[54],c49[55],s49[54]);


full_add fa49_55(s48[56],c48[56],andpr51[55],c49[56],s49[55]);


full_add fa49_56(s48[57],c48[57],andpr51[56],c49[57],s49[56]);


full_add fa49_57(s48[58],c48[58],andpr51[57],c49[58],s49[57]);


full_add fa49_58(s48[59],c48[59],andpr51[58],c49[59],s49[58]);


full_add fa49_59(s48[60],c48[60],andpr51[59],c49[60],s49[59]);


full_add fa49_60(s48[61],c48[61],andpr51[60],c49[61],s49[60]);


full_add fa49_61(s48[62],c48[62],andpr51[61],c49[62],s49[61]);


full_add fa49_62(si[49],c48[63],andpr51[62],c49[63],s49[62]);



half_adder ha50(s49[0],c49[0],c50[0],p[50]);


full_add fa50_0(s49[1],c49[1],andpr52[0],c50[1],s50[0]);


full_add fa50_1(s49[2],c49[2],andpr52[1],c50[2],s50[1]);


full_add fa50_2(s49[3],c49[3],andpr52[2],c50[3],s50[2]);


full_add fa50_3(s49[4],c49[4],andpr52[3],c50[4],s50[3]);


full_add fa50_4(s49[5],c49[5],andpr52[4],c50[5],s50[4]);


full_add fa50_5(s49[6],c49[6],andpr52[5],c50[6],s50[5]);


full_add fa50_6(s49[7],c49[7],andpr52[6],c50[7],s50[6]);


full_add fa50_7(s49[8],c49[8],andpr52[7],c50[8],s50[7]);


full_add fa50_8(s49[9],c49[9],andpr52[8],c50[9],s50[8]);


full_add fa50_9(s49[10],c49[10],andpr52[9],c50[10],s50[9]);


full_add fa50_10(s49[11],c49[11],andpr52[10],c50[11],s50[10]);


full_add fa50_11(s49[12],c49[12],andpr52[11],c50[12],s50[11]);


full_add fa50_12(s49[13],c49[13],andpr52[12],c50[13],s50[12]);


full_add fa50_13(s49[14],c49[14],andpr52[13],c50[14],s50[13]);


full_add fa50_14(s49[15],c49[15],andpr52[14],c50[15],s50[14]);


full_add fa50_15(s49[16],c49[16],andpr52[15],c50[16],s50[15]);


full_add fa50_16(s49[17],c49[17],andpr52[16],c50[17],s50[16]);


full_add fa50_17(s49[18],c49[18],andpr52[17],c50[18],s50[17]);


full_add fa50_18(s49[19],c49[19],andpr52[18],c50[19],s50[18]);


full_add fa50_19(s49[20],c49[20],andpr52[19],c50[20],s50[19]);


full_add fa50_20(s49[21],c49[21],andpr52[20],c50[21],s50[20]);


full_add fa50_21(s49[22],c49[22],andpr52[21],c50[22],s50[21]);


full_add fa50_22(s49[23],c49[23],andpr52[22],c50[23],s50[22]);


full_add fa50_23(s49[24],c49[24],andpr52[23],c50[24],s50[23]);


full_add fa50_24(s49[25],c49[25],andpr52[24],c50[25],s50[24]);


full_add fa50_25(s49[26],c49[26],andpr52[25],c50[26],s50[25]);


full_add fa50_26(s49[27],c49[27],andpr52[26],c50[27],s50[26]);


full_add fa50_27(s49[28],c49[28],andpr52[27],c50[28],s50[27]);


full_add fa50_28(s49[29],c49[29],andpr52[28],c50[29],s50[28]);


full_add fa50_29(s49[30],c49[30],andpr52[29],c50[30],s50[29]);


full_add fa50_30(s49[31],c49[31],andpr52[30],c50[31],s50[30]);


full_add fa50_31(s49[32],c49[32],andpr52[31],c50[32],s50[31]);


full_add fa50_32(s49[33],c49[33],andpr52[32],c50[33],s50[32]);


full_add fa50_33(s49[34],c49[34],andpr52[33],c50[34],s50[33]);


full_add fa50_34(s49[35],c49[35],andpr52[34],c50[35],s50[34]);


full_add fa50_35(s49[36],c49[36],andpr52[35],c50[36],s50[35]);


full_add fa50_36(s49[37],c49[37],andpr52[36],c50[37],s50[36]);


full_add fa50_37(s49[38],c49[38],andpr52[37],c50[38],s50[37]);


full_add fa50_38(s49[39],c49[39],andpr52[38],c50[39],s50[38]);


full_add fa50_39(s49[40],c49[40],andpr52[39],c50[40],s50[39]);


full_add fa50_40(s49[41],c49[41],andpr52[40],c50[41],s50[40]);


full_add fa50_41(s49[42],c49[42],andpr52[41],c50[42],s50[41]);


full_add fa50_42(s49[43],c49[43],andpr52[42],c50[43],s50[42]);


full_add fa50_43(s49[44],c49[44],andpr52[43],c50[44],s50[43]);


full_add fa50_44(s49[45],c49[45],andpr52[44],c50[45],s50[44]);


full_add fa50_45(s49[46],c49[46],andpr52[45],c50[46],s50[45]);


full_add fa50_46(s49[47],c49[47],andpr52[46],c50[47],s50[46]);


full_add fa50_47(s49[48],c49[48],andpr52[47],c50[48],s50[47]);


full_add fa50_48(s49[49],c49[49],andpr52[48],c50[49],s50[48]);


full_add fa50_49(s49[50],c49[50],andpr52[49],c50[50],s50[49]);


full_add fa50_50(s49[51],c49[51],andpr52[50],c50[51],s50[50]);


full_add fa50_51(s49[52],c49[52],andpr52[51],c50[52],s50[51]);


full_add fa50_52(s49[53],c49[53],andpr52[52],c50[53],s50[52]);


full_add fa50_53(s49[54],c49[54],andpr52[53],c50[54],s50[53]);


full_add fa50_54(s49[55],c49[55],andpr52[54],c50[55],s50[54]);


full_add fa50_55(s49[56],c49[56],andpr52[55],c50[56],s50[55]);


full_add fa50_56(s49[57],c49[57],andpr52[56],c50[57],s50[56]);


full_add fa50_57(s49[58],c49[58],andpr52[57],c50[58],s50[57]);


full_add fa50_58(s49[59],c49[59],andpr52[58],c50[59],s50[58]);


full_add fa50_59(s49[60],c49[60],andpr52[59],c50[60],s50[59]);


full_add fa50_60(s49[61],c49[61],andpr52[60],c50[61],s50[60]);


full_add fa50_61(s49[62],c49[62],andpr52[61],c50[62],s50[61]);


full_add fa50_62(si[50],c49[63],andpr52[62],c50[63],s50[62]);



half_adder ha51(s50[0],c50[0],c51[0],p[51]);


full_add fa51_0(s50[1],c50[1],andpr53[0],c51[1],s51[0]);


full_add fa51_1(s50[2],c50[2],andpr53[1],c51[2],s51[1]);


full_add fa51_2(s50[3],c50[3],andpr53[2],c51[3],s51[2]);


full_add fa51_3(s50[4],c50[4],andpr53[3],c51[4],s51[3]);


full_add fa51_4(s50[5],c50[5],andpr53[4],c51[5],s51[4]);


full_add fa51_5(s50[6],c50[6],andpr53[5],c51[6],s51[5]);


full_add fa51_6(s50[7],c50[7],andpr53[6],c51[7],s51[6]);


full_add fa51_7(s50[8],c50[8],andpr53[7],c51[8],s51[7]);


full_add fa51_8(s50[9],c50[9],andpr53[8],c51[9],s51[8]);


full_add fa51_9(s50[10],c50[10],andpr53[9],c51[10],s51[9]);


full_add fa51_10(s50[11],c50[11],andpr53[10],c51[11],s51[10]);


full_add fa51_11(s50[12],c50[12],andpr53[11],c51[12],s51[11]);


full_add fa51_12(s50[13],c50[13],andpr53[12],c51[13],s51[12]);


full_add fa51_13(s50[14],c50[14],andpr53[13],c51[14],s51[13]);


full_add fa51_14(s50[15],c50[15],andpr53[14],c51[15],s51[14]);


full_add fa51_15(s50[16],c50[16],andpr53[15],c51[16],s51[15]);


full_add fa51_16(s50[17],c50[17],andpr53[16],c51[17],s51[16]);


full_add fa51_17(s50[18],c50[18],andpr53[17],c51[18],s51[17]);


full_add fa51_18(s50[19],c50[19],andpr53[18],c51[19],s51[18]);


full_add fa51_19(s50[20],c50[20],andpr53[19],c51[20],s51[19]);


full_add fa51_20(s50[21],c50[21],andpr53[20],c51[21],s51[20]);


full_add fa51_21(s50[22],c50[22],andpr53[21],c51[22],s51[21]);


full_add fa51_22(s50[23],c50[23],andpr53[22],c51[23],s51[22]);


full_add fa51_23(s50[24],c50[24],andpr53[23],c51[24],s51[23]);


full_add fa51_24(s50[25],c50[25],andpr53[24],c51[25],s51[24]);


full_add fa51_25(s50[26],c50[26],andpr53[25],c51[26],s51[25]);


full_add fa51_26(s50[27],c50[27],andpr53[26],c51[27],s51[26]);


full_add fa51_27(s50[28],c50[28],andpr53[27],c51[28],s51[27]);


full_add fa51_28(s50[29],c50[29],andpr53[28],c51[29],s51[28]);


full_add fa51_29(s50[30],c50[30],andpr53[29],c51[30],s51[29]);


full_add fa51_30(s50[31],c50[31],andpr53[30],c51[31],s51[30]);


full_add fa51_31(s50[32],c50[32],andpr53[31],c51[32],s51[31]);


full_add fa51_32(s50[33],c50[33],andpr53[32],c51[33],s51[32]);


full_add fa51_33(s50[34],c50[34],andpr53[33],c51[34],s51[33]);


full_add fa51_34(s50[35],c50[35],andpr53[34],c51[35],s51[34]);


full_add fa51_35(s50[36],c50[36],andpr53[35],c51[36],s51[35]);


full_add fa51_36(s50[37],c50[37],andpr53[36],c51[37],s51[36]);


full_add fa51_37(s50[38],c50[38],andpr53[37],c51[38],s51[37]);


full_add fa51_38(s50[39],c50[39],andpr53[38],c51[39],s51[38]);


full_add fa51_39(s50[40],c50[40],andpr53[39],c51[40],s51[39]);


full_add fa51_40(s50[41],c50[41],andpr53[40],c51[41],s51[40]);


full_add fa51_41(s50[42],c50[42],andpr53[41],c51[42],s51[41]);


full_add fa51_42(s50[43],c50[43],andpr53[42],c51[43],s51[42]);


full_add fa51_43(s50[44],c50[44],andpr53[43],c51[44],s51[43]);


full_add fa51_44(s50[45],c50[45],andpr53[44],c51[45],s51[44]);


full_add fa51_45(s50[46],c50[46],andpr53[45],c51[46],s51[45]);


full_add fa51_46(s50[47],c50[47],andpr53[46],c51[47],s51[46]);


full_add fa51_47(s50[48],c50[48],andpr53[47],c51[48],s51[47]);


full_add fa51_48(s50[49],c50[49],andpr53[48],c51[49],s51[48]);


full_add fa51_49(s50[50],c50[50],andpr53[49],c51[50],s51[49]);


full_add fa51_50(s50[51],c50[51],andpr53[50],c51[51],s51[50]);


full_add fa51_51(s50[52],c50[52],andpr53[51],c51[52],s51[51]);


full_add fa51_52(s50[53],c50[53],andpr53[52],c51[53],s51[52]);


full_add fa51_53(s50[54],c50[54],andpr53[53],c51[54],s51[53]);


full_add fa51_54(s50[55],c50[55],andpr53[54],c51[55],s51[54]);


full_add fa51_55(s50[56],c50[56],andpr53[55],c51[56],s51[55]);


full_add fa51_56(s50[57],c50[57],andpr53[56],c51[57],s51[56]);


full_add fa51_57(s50[58],c50[58],andpr53[57],c51[58],s51[57]);


full_add fa51_58(s50[59],c50[59],andpr53[58],c51[59],s51[58]);


full_add fa51_59(s50[60],c50[60],andpr53[59],c51[60],s51[59]);


full_add fa51_60(s50[61],c50[61],andpr53[60],c51[61],s51[60]);


full_add fa51_61(s50[62],c50[62],andpr53[61],c51[62],s51[61]);


full_add fa51_62(si[51],c50[63],andpr53[62],c51[63],s51[62]);



half_adder ha52(s51[0],c51[0],c52[0],p[52]);


full_add fa52_0(s51[1],c51[1],andpr54[0],c52[1],s52[0]);


full_add fa52_1(s51[2],c51[2],andpr54[1],c52[2],s52[1]);


full_add fa52_2(s51[3],c51[3],andpr54[2],c52[3],s52[2]);


full_add fa52_3(s51[4],c51[4],andpr54[3],c52[4],s52[3]);


full_add fa52_4(s51[5],c51[5],andpr54[4],c52[5],s52[4]);


full_add fa52_5(s51[6],c51[6],andpr54[5],c52[6],s52[5]);


full_add fa52_6(s51[7],c51[7],andpr54[6],c52[7],s52[6]);


full_add fa52_7(s51[8],c51[8],andpr54[7],c52[8],s52[7]);


full_add fa52_8(s51[9],c51[9],andpr54[8],c52[9],s52[8]);


full_add fa52_9(s51[10],c51[10],andpr54[9],c52[10],s52[9]);


full_add fa52_10(s51[11],c51[11],andpr54[10],c52[11],s52[10]);


full_add fa52_11(s51[12],c51[12],andpr54[11],c52[12],s52[11]);


full_add fa52_12(s51[13],c51[13],andpr54[12],c52[13],s52[12]);


full_add fa52_13(s51[14],c51[14],andpr54[13],c52[14],s52[13]);


full_add fa52_14(s51[15],c51[15],andpr54[14],c52[15],s52[14]);


full_add fa52_15(s51[16],c51[16],andpr54[15],c52[16],s52[15]);


full_add fa52_16(s51[17],c51[17],andpr54[16],c52[17],s52[16]);


full_add fa52_17(s51[18],c51[18],andpr54[17],c52[18],s52[17]);


full_add fa52_18(s51[19],c51[19],andpr54[18],c52[19],s52[18]);


full_add fa52_19(s51[20],c51[20],andpr54[19],c52[20],s52[19]);


full_add fa52_20(s51[21],c51[21],andpr54[20],c52[21],s52[20]);


full_add fa52_21(s51[22],c51[22],andpr54[21],c52[22],s52[21]);


full_add fa52_22(s51[23],c51[23],andpr54[22],c52[23],s52[22]);


full_add fa52_23(s51[24],c51[24],andpr54[23],c52[24],s52[23]);


full_add fa52_24(s51[25],c51[25],andpr54[24],c52[25],s52[24]);


full_add fa52_25(s51[26],c51[26],andpr54[25],c52[26],s52[25]);


full_add fa52_26(s51[27],c51[27],andpr54[26],c52[27],s52[26]);


full_add fa52_27(s51[28],c51[28],andpr54[27],c52[28],s52[27]);


full_add fa52_28(s51[29],c51[29],andpr54[28],c52[29],s52[28]);


full_add fa52_29(s51[30],c51[30],andpr54[29],c52[30],s52[29]);


full_add fa52_30(s51[31],c51[31],andpr54[30],c52[31],s52[30]);


full_add fa52_31(s51[32],c51[32],andpr54[31],c52[32],s52[31]);


full_add fa52_32(s51[33],c51[33],andpr54[32],c52[33],s52[32]);


full_add fa52_33(s51[34],c51[34],andpr54[33],c52[34],s52[33]);


full_add fa52_34(s51[35],c51[35],andpr54[34],c52[35],s52[34]);


full_add fa52_35(s51[36],c51[36],andpr54[35],c52[36],s52[35]);


full_add fa52_36(s51[37],c51[37],andpr54[36],c52[37],s52[36]);


full_add fa52_37(s51[38],c51[38],andpr54[37],c52[38],s52[37]);


full_add fa52_38(s51[39],c51[39],andpr54[38],c52[39],s52[38]);


full_add fa52_39(s51[40],c51[40],andpr54[39],c52[40],s52[39]);


full_add fa52_40(s51[41],c51[41],andpr54[40],c52[41],s52[40]);


full_add fa52_41(s51[42],c51[42],andpr54[41],c52[42],s52[41]);


full_add fa52_42(s51[43],c51[43],andpr54[42],c52[43],s52[42]);


full_add fa52_43(s51[44],c51[44],andpr54[43],c52[44],s52[43]);


full_add fa52_44(s51[45],c51[45],andpr54[44],c52[45],s52[44]);


full_add fa52_45(s51[46],c51[46],andpr54[45],c52[46],s52[45]);


full_add fa52_46(s51[47],c51[47],andpr54[46],c52[47],s52[46]);


full_add fa52_47(s51[48],c51[48],andpr54[47],c52[48],s52[47]);


full_add fa52_48(s51[49],c51[49],andpr54[48],c52[49],s52[48]);


full_add fa52_49(s51[50],c51[50],andpr54[49],c52[50],s52[49]);


full_add fa52_50(s51[51],c51[51],andpr54[50],c52[51],s52[50]);


full_add fa52_51(s51[52],c51[52],andpr54[51],c52[52],s52[51]);


full_add fa52_52(s51[53],c51[53],andpr54[52],c52[53],s52[52]);


full_add fa52_53(s51[54],c51[54],andpr54[53],c52[54],s52[53]);


full_add fa52_54(s51[55],c51[55],andpr54[54],c52[55],s52[54]);


full_add fa52_55(s51[56],c51[56],andpr54[55],c52[56],s52[55]);


full_add fa52_56(s51[57],c51[57],andpr54[56],c52[57],s52[56]);


full_add fa52_57(s51[58],c51[58],andpr54[57],c52[58],s52[57]);


full_add fa52_58(s51[59],c51[59],andpr54[58],c52[59],s52[58]);


full_add fa52_59(s51[60],c51[60],andpr54[59],c52[60],s52[59]);


full_add fa52_60(s51[61],c51[61],andpr54[60],c52[61],s52[60]);


full_add fa52_61(s51[62],c51[62],andpr54[61],c52[62],s52[61]);


full_add fa52_62(si[52],c51[63],andpr54[62],c52[63],s52[62]);



half_adder ha53(s52[0],c52[0],c53[0],p[53]);


full_add fa53_0(s52[1],c52[1],andpr55[0],c53[1],s53[0]);


full_add fa53_1(s52[2],c52[2],andpr55[1],c53[2],s53[1]);


full_add fa53_2(s52[3],c52[3],andpr55[2],c53[3],s53[2]);


full_add fa53_3(s52[4],c52[4],andpr55[3],c53[4],s53[3]);


full_add fa53_4(s52[5],c52[5],andpr55[4],c53[5],s53[4]);


full_add fa53_5(s52[6],c52[6],andpr55[5],c53[6],s53[5]);


full_add fa53_6(s52[7],c52[7],andpr55[6],c53[7],s53[6]);


full_add fa53_7(s52[8],c52[8],andpr55[7],c53[8],s53[7]);


full_add fa53_8(s52[9],c52[9],andpr55[8],c53[9],s53[8]);


full_add fa53_9(s52[10],c52[10],andpr55[9],c53[10],s53[9]);


full_add fa53_10(s52[11],c52[11],andpr55[10],c53[11],s53[10]);


full_add fa53_11(s52[12],c52[12],andpr55[11],c53[12],s53[11]);


full_add fa53_12(s52[13],c52[13],andpr55[12],c53[13],s53[12]);


full_add fa53_13(s52[14],c52[14],andpr55[13],c53[14],s53[13]);


full_add fa53_14(s52[15],c52[15],andpr55[14],c53[15],s53[14]);


full_add fa53_15(s52[16],c52[16],andpr55[15],c53[16],s53[15]);


full_add fa53_16(s52[17],c52[17],andpr55[16],c53[17],s53[16]);


full_add fa53_17(s52[18],c52[18],andpr55[17],c53[18],s53[17]);


full_add fa53_18(s52[19],c52[19],andpr55[18],c53[19],s53[18]);


full_add fa53_19(s52[20],c52[20],andpr55[19],c53[20],s53[19]);


full_add fa53_20(s52[21],c52[21],andpr55[20],c53[21],s53[20]);


full_add fa53_21(s52[22],c52[22],andpr55[21],c53[22],s53[21]);


full_add fa53_22(s52[23],c52[23],andpr55[22],c53[23],s53[22]);


full_add fa53_23(s52[24],c52[24],andpr55[23],c53[24],s53[23]);


full_add fa53_24(s52[25],c52[25],andpr55[24],c53[25],s53[24]);


full_add fa53_25(s52[26],c52[26],andpr55[25],c53[26],s53[25]);


full_add fa53_26(s52[27],c52[27],andpr55[26],c53[27],s53[26]);


full_add fa53_27(s52[28],c52[28],andpr55[27],c53[28],s53[27]);


full_add fa53_28(s52[29],c52[29],andpr55[28],c53[29],s53[28]);


full_add fa53_29(s52[30],c52[30],andpr55[29],c53[30],s53[29]);


full_add fa53_30(s52[31],c52[31],andpr55[30],c53[31],s53[30]);


full_add fa53_31(s52[32],c52[32],andpr55[31],c53[32],s53[31]);


full_add fa53_32(s52[33],c52[33],andpr55[32],c53[33],s53[32]);


full_add fa53_33(s52[34],c52[34],andpr55[33],c53[34],s53[33]);


full_add fa53_34(s52[35],c52[35],andpr55[34],c53[35],s53[34]);


full_add fa53_35(s52[36],c52[36],andpr55[35],c53[36],s53[35]);


full_add fa53_36(s52[37],c52[37],andpr55[36],c53[37],s53[36]);


full_add fa53_37(s52[38],c52[38],andpr55[37],c53[38],s53[37]);


full_add fa53_38(s52[39],c52[39],andpr55[38],c53[39],s53[38]);


full_add fa53_39(s52[40],c52[40],andpr55[39],c53[40],s53[39]);


full_add fa53_40(s52[41],c52[41],andpr55[40],c53[41],s53[40]);


full_add fa53_41(s52[42],c52[42],andpr55[41],c53[42],s53[41]);


full_add fa53_42(s52[43],c52[43],andpr55[42],c53[43],s53[42]);


full_add fa53_43(s52[44],c52[44],andpr55[43],c53[44],s53[43]);


full_add fa53_44(s52[45],c52[45],andpr55[44],c53[45],s53[44]);


full_add fa53_45(s52[46],c52[46],andpr55[45],c53[46],s53[45]);


full_add fa53_46(s52[47],c52[47],andpr55[46],c53[47],s53[46]);


full_add fa53_47(s52[48],c52[48],andpr55[47],c53[48],s53[47]);


full_add fa53_48(s52[49],c52[49],andpr55[48],c53[49],s53[48]);


full_add fa53_49(s52[50],c52[50],andpr55[49],c53[50],s53[49]);


full_add fa53_50(s52[51],c52[51],andpr55[50],c53[51],s53[50]);


full_add fa53_51(s52[52],c52[52],andpr55[51],c53[52],s53[51]);


full_add fa53_52(s52[53],c52[53],andpr55[52],c53[53],s53[52]);


full_add fa53_53(s52[54],c52[54],andpr55[53],c53[54],s53[53]);


full_add fa53_54(s52[55],c52[55],andpr55[54],c53[55],s53[54]);


full_add fa53_55(s52[56],c52[56],andpr55[55],c53[56],s53[55]);


full_add fa53_56(s52[57],c52[57],andpr55[56],c53[57],s53[56]);


full_add fa53_57(s52[58],c52[58],andpr55[57],c53[58],s53[57]);


full_add fa53_58(s52[59],c52[59],andpr55[58],c53[59],s53[58]);


full_add fa53_59(s52[60],c52[60],andpr55[59],c53[60],s53[59]);


full_add fa53_60(s52[61],c52[61],andpr55[60],c53[61],s53[60]);


full_add fa53_61(s52[62],c52[62],andpr55[61],c53[62],s53[61]);


full_add fa53_62(si[53],c52[63],andpr55[62],c53[63],s53[62]);



half_adder ha54(s53[0],c53[0],c54[0],p[54]);


full_add fa54_0(s53[1],c53[1],andpr56[0],c54[1],s54[0]);


full_add fa54_1(s53[2],c53[2],andpr56[1],c54[2],s54[1]);


full_add fa54_2(s53[3],c53[3],andpr56[2],c54[3],s54[2]);


full_add fa54_3(s53[4],c53[4],andpr56[3],c54[4],s54[3]);


full_add fa54_4(s53[5],c53[5],andpr56[4],c54[5],s54[4]);


full_add fa54_5(s53[6],c53[6],andpr56[5],c54[6],s54[5]);


full_add fa54_6(s53[7],c53[7],andpr56[6],c54[7],s54[6]);


full_add fa54_7(s53[8],c53[8],andpr56[7],c54[8],s54[7]);


full_add fa54_8(s53[9],c53[9],andpr56[8],c54[9],s54[8]);


full_add fa54_9(s53[10],c53[10],andpr56[9],c54[10],s54[9]);


full_add fa54_10(s53[11],c53[11],andpr56[10],c54[11],s54[10]);


full_add fa54_11(s53[12],c53[12],andpr56[11],c54[12],s54[11]);


full_add fa54_12(s53[13],c53[13],andpr56[12],c54[13],s54[12]);


full_add fa54_13(s53[14],c53[14],andpr56[13],c54[14],s54[13]);


full_add fa54_14(s53[15],c53[15],andpr56[14],c54[15],s54[14]);


full_add fa54_15(s53[16],c53[16],andpr56[15],c54[16],s54[15]);


full_add fa54_16(s53[17],c53[17],andpr56[16],c54[17],s54[16]);


full_add fa54_17(s53[18],c53[18],andpr56[17],c54[18],s54[17]);


full_add fa54_18(s53[19],c53[19],andpr56[18],c54[19],s54[18]);


full_add fa54_19(s53[20],c53[20],andpr56[19],c54[20],s54[19]);


full_add fa54_20(s53[21],c53[21],andpr56[20],c54[21],s54[20]);


full_add fa54_21(s53[22],c53[22],andpr56[21],c54[22],s54[21]);


full_add fa54_22(s53[23],c53[23],andpr56[22],c54[23],s54[22]);


full_add fa54_23(s53[24],c53[24],andpr56[23],c54[24],s54[23]);


full_add fa54_24(s53[25],c53[25],andpr56[24],c54[25],s54[24]);


full_add fa54_25(s53[26],c53[26],andpr56[25],c54[26],s54[25]);


full_add fa54_26(s53[27],c53[27],andpr56[26],c54[27],s54[26]);


full_add fa54_27(s53[28],c53[28],andpr56[27],c54[28],s54[27]);


full_add fa54_28(s53[29],c53[29],andpr56[28],c54[29],s54[28]);


full_add fa54_29(s53[30],c53[30],andpr56[29],c54[30],s54[29]);


full_add fa54_30(s53[31],c53[31],andpr56[30],c54[31],s54[30]);


full_add fa54_31(s53[32],c53[32],andpr56[31],c54[32],s54[31]);


full_add fa54_32(s53[33],c53[33],andpr56[32],c54[33],s54[32]);


full_add fa54_33(s53[34],c53[34],andpr56[33],c54[34],s54[33]);


full_add fa54_34(s53[35],c53[35],andpr56[34],c54[35],s54[34]);


full_add fa54_35(s53[36],c53[36],andpr56[35],c54[36],s54[35]);


full_add fa54_36(s53[37],c53[37],andpr56[36],c54[37],s54[36]);


full_add fa54_37(s53[38],c53[38],andpr56[37],c54[38],s54[37]);


full_add fa54_38(s53[39],c53[39],andpr56[38],c54[39],s54[38]);


full_add fa54_39(s53[40],c53[40],andpr56[39],c54[40],s54[39]);


full_add fa54_40(s53[41],c53[41],andpr56[40],c54[41],s54[40]);


full_add fa54_41(s53[42],c53[42],andpr56[41],c54[42],s54[41]);


full_add fa54_42(s53[43],c53[43],andpr56[42],c54[43],s54[42]);


full_add fa54_43(s53[44],c53[44],andpr56[43],c54[44],s54[43]);


full_add fa54_44(s53[45],c53[45],andpr56[44],c54[45],s54[44]);


full_add fa54_45(s53[46],c53[46],andpr56[45],c54[46],s54[45]);


full_add fa54_46(s53[47],c53[47],andpr56[46],c54[47],s54[46]);


full_add fa54_47(s53[48],c53[48],andpr56[47],c54[48],s54[47]);


full_add fa54_48(s53[49],c53[49],andpr56[48],c54[49],s54[48]);


full_add fa54_49(s53[50],c53[50],andpr56[49],c54[50],s54[49]);


full_add fa54_50(s53[51],c53[51],andpr56[50],c54[51],s54[50]);


full_add fa54_51(s53[52],c53[52],andpr56[51],c54[52],s54[51]);


full_add fa54_52(s53[53],c53[53],andpr56[52],c54[53],s54[52]);


full_add fa54_53(s53[54],c53[54],andpr56[53],c54[54],s54[53]);


full_add fa54_54(s53[55],c53[55],andpr56[54],c54[55],s54[54]);


full_add fa54_55(s53[56],c53[56],andpr56[55],c54[56],s54[55]);


full_add fa54_56(s53[57],c53[57],andpr56[56],c54[57],s54[56]);


full_add fa54_57(s53[58],c53[58],andpr56[57],c54[58],s54[57]);


full_add fa54_58(s53[59],c53[59],andpr56[58],c54[59],s54[58]);


full_add fa54_59(s53[60],c53[60],andpr56[59],c54[60],s54[59]);


full_add fa54_60(s53[61],c53[61],andpr56[60],c54[61],s54[60]);


full_add fa54_61(s53[62],c53[62],andpr56[61],c54[62],s54[61]);


full_add fa54_62(si[54],c53[63],andpr56[62],c54[63],s54[62]);



half_adder ha55(s54[0],c54[0],c55[0],p[55]);


full_add fa55_0(s54[1],c54[1],andpr57[0],c55[1],s55[0]);


full_add fa55_1(s54[2],c54[2],andpr57[1],c55[2],s55[1]);


full_add fa55_2(s54[3],c54[3],andpr57[2],c55[3],s55[2]);


full_add fa55_3(s54[4],c54[4],andpr57[3],c55[4],s55[3]);


full_add fa55_4(s54[5],c54[5],andpr57[4],c55[5],s55[4]);


full_add fa55_5(s54[6],c54[6],andpr57[5],c55[6],s55[5]);


full_add fa55_6(s54[7],c54[7],andpr57[6],c55[7],s55[6]);


full_add fa55_7(s54[8],c54[8],andpr57[7],c55[8],s55[7]);


full_add fa55_8(s54[9],c54[9],andpr57[8],c55[9],s55[8]);


full_add fa55_9(s54[10],c54[10],andpr57[9],c55[10],s55[9]);


full_add fa55_10(s54[11],c54[11],andpr57[10],c55[11],s55[10]);


full_add fa55_11(s54[12],c54[12],andpr57[11],c55[12],s55[11]);


full_add fa55_12(s54[13],c54[13],andpr57[12],c55[13],s55[12]);


full_add fa55_13(s54[14],c54[14],andpr57[13],c55[14],s55[13]);


full_add fa55_14(s54[15],c54[15],andpr57[14],c55[15],s55[14]);


full_add fa55_15(s54[16],c54[16],andpr57[15],c55[16],s55[15]);


full_add fa55_16(s54[17],c54[17],andpr57[16],c55[17],s55[16]);


full_add fa55_17(s54[18],c54[18],andpr57[17],c55[18],s55[17]);


full_add fa55_18(s54[19],c54[19],andpr57[18],c55[19],s55[18]);


full_add fa55_19(s54[20],c54[20],andpr57[19],c55[20],s55[19]);


full_add fa55_20(s54[21],c54[21],andpr57[20],c55[21],s55[20]);


full_add fa55_21(s54[22],c54[22],andpr57[21],c55[22],s55[21]);


full_add fa55_22(s54[23],c54[23],andpr57[22],c55[23],s55[22]);


full_add fa55_23(s54[24],c54[24],andpr57[23],c55[24],s55[23]);


full_add fa55_24(s54[25],c54[25],andpr57[24],c55[25],s55[24]);


full_add fa55_25(s54[26],c54[26],andpr57[25],c55[26],s55[25]);


full_add fa55_26(s54[27],c54[27],andpr57[26],c55[27],s55[26]);


full_add fa55_27(s54[28],c54[28],andpr57[27],c55[28],s55[27]);


full_add fa55_28(s54[29],c54[29],andpr57[28],c55[29],s55[28]);


full_add fa55_29(s54[30],c54[30],andpr57[29],c55[30],s55[29]);


full_add fa55_30(s54[31],c54[31],andpr57[30],c55[31],s55[30]);


full_add fa55_31(s54[32],c54[32],andpr57[31],c55[32],s55[31]);


full_add fa55_32(s54[33],c54[33],andpr57[32],c55[33],s55[32]);


full_add fa55_33(s54[34],c54[34],andpr57[33],c55[34],s55[33]);


full_add fa55_34(s54[35],c54[35],andpr57[34],c55[35],s55[34]);


full_add fa55_35(s54[36],c54[36],andpr57[35],c55[36],s55[35]);


full_add fa55_36(s54[37],c54[37],andpr57[36],c55[37],s55[36]);


full_add fa55_37(s54[38],c54[38],andpr57[37],c55[38],s55[37]);


full_add fa55_38(s54[39],c54[39],andpr57[38],c55[39],s55[38]);


full_add fa55_39(s54[40],c54[40],andpr57[39],c55[40],s55[39]);


full_add fa55_40(s54[41],c54[41],andpr57[40],c55[41],s55[40]);


full_add fa55_41(s54[42],c54[42],andpr57[41],c55[42],s55[41]);


full_add fa55_42(s54[43],c54[43],andpr57[42],c55[43],s55[42]);


full_add fa55_43(s54[44],c54[44],andpr57[43],c55[44],s55[43]);


full_add fa55_44(s54[45],c54[45],andpr57[44],c55[45],s55[44]);


full_add fa55_45(s54[46],c54[46],andpr57[45],c55[46],s55[45]);


full_add fa55_46(s54[47],c54[47],andpr57[46],c55[47],s55[46]);


full_add fa55_47(s54[48],c54[48],andpr57[47],c55[48],s55[47]);


full_add fa55_48(s54[49],c54[49],andpr57[48],c55[49],s55[48]);


full_add fa55_49(s54[50],c54[50],andpr57[49],c55[50],s55[49]);


full_add fa55_50(s54[51],c54[51],andpr57[50],c55[51],s55[50]);


full_add fa55_51(s54[52],c54[52],andpr57[51],c55[52],s55[51]);


full_add fa55_52(s54[53],c54[53],andpr57[52],c55[53],s55[52]);


full_add fa55_53(s54[54],c54[54],andpr57[53],c55[54],s55[53]);


full_add fa55_54(s54[55],c54[55],andpr57[54],c55[55],s55[54]);


full_add fa55_55(s54[56],c54[56],andpr57[55],c55[56],s55[55]);


full_add fa55_56(s54[57],c54[57],andpr57[56],c55[57],s55[56]);


full_add fa55_57(s54[58],c54[58],andpr57[57],c55[58],s55[57]);


full_add fa55_58(s54[59],c54[59],andpr57[58],c55[59],s55[58]);


full_add fa55_59(s54[60],c54[60],andpr57[59],c55[60],s55[59]);


full_add fa55_60(s54[61],c54[61],andpr57[60],c55[61],s55[60]);


full_add fa55_61(s54[62],c54[62],andpr57[61],c55[62],s55[61]);


full_add fa55_62(si[55],c54[63],andpr57[62],c55[63],s55[62]);



half_adder ha56(s55[0],c55[0],c56[0],p[56]);


full_add fa56_0(s55[1],c55[1],andpr58[0],c56[1],s56[0]);


full_add fa56_1(s55[2],c55[2],andpr58[1],c56[2],s56[1]);


full_add fa56_2(s55[3],c55[3],andpr58[2],c56[3],s56[2]);


full_add fa56_3(s55[4],c55[4],andpr58[3],c56[4],s56[3]);


full_add fa56_4(s55[5],c55[5],andpr58[4],c56[5],s56[4]);


full_add fa56_5(s55[6],c55[6],andpr58[5],c56[6],s56[5]);


full_add fa56_6(s55[7],c55[7],andpr58[6],c56[7],s56[6]);


full_add fa56_7(s55[8],c55[8],andpr58[7],c56[8],s56[7]);


full_add fa56_8(s55[9],c55[9],andpr58[8],c56[9],s56[8]);


full_add fa56_9(s55[10],c55[10],andpr58[9],c56[10],s56[9]);


full_add fa56_10(s55[11],c55[11],andpr58[10],c56[11],s56[10]);


full_add fa56_11(s55[12],c55[12],andpr58[11],c56[12],s56[11]);


full_add fa56_12(s55[13],c55[13],andpr58[12],c56[13],s56[12]);


full_add fa56_13(s55[14],c55[14],andpr58[13],c56[14],s56[13]);


full_add fa56_14(s55[15],c55[15],andpr58[14],c56[15],s56[14]);


full_add fa56_15(s55[16],c55[16],andpr58[15],c56[16],s56[15]);


full_add fa56_16(s55[17],c55[17],andpr58[16],c56[17],s56[16]);


full_add fa56_17(s55[18],c55[18],andpr58[17],c56[18],s56[17]);


full_add fa56_18(s55[19],c55[19],andpr58[18],c56[19],s56[18]);


full_add fa56_19(s55[20],c55[20],andpr58[19],c56[20],s56[19]);


full_add fa56_20(s55[21],c55[21],andpr58[20],c56[21],s56[20]);


full_add fa56_21(s55[22],c55[22],andpr58[21],c56[22],s56[21]);


full_add fa56_22(s55[23],c55[23],andpr58[22],c56[23],s56[22]);


full_add fa56_23(s55[24],c55[24],andpr58[23],c56[24],s56[23]);


full_add fa56_24(s55[25],c55[25],andpr58[24],c56[25],s56[24]);


full_add fa56_25(s55[26],c55[26],andpr58[25],c56[26],s56[25]);


full_add fa56_26(s55[27],c55[27],andpr58[26],c56[27],s56[26]);


full_add fa56_27(s55[28],c55[28],andpr58[27],c56[28],s56[27]);


full_add fa56_28(s55[29],c55[29],andpr58[28],c56[29],s56[28]);


full_add fa56_29(s55[30],c55[30],andpr58[29],c56[30],s56[29]);


full_add fa56_30(s55[31],c55[31],andpr58[30],c56[31],s56[30]);


full_add fa56_31(s55[32],c55[32],andpr58[31],c56[32],s56[31]);


full_add fa56_32(s55[33],c55[33],andpr58[32],c56[33],s56[32]);


full_add fa56_33(s55[34],c55[34],andpr58[33],c56[34],s56[33]);


full_add fa56_34(s55[35],c55[35],andpr58[34],c56[35],s56[34]);


full_add fa56_35(s55[36],c55[36],andpr58[35],c56[36],s56[35]);


full_add fa56_36(s55[37],c55[37],andpr58[36],c56[37],s56[36]);


full_add fa56_37(s55[38],c55[38],andpr58[37],c56[38],s56[37]);


full_add fa56_38(s55[39],c55[39],andpr58[38],c56[39],s56[38]);


full_add fa56_39(s55[40],c55[40],andpr58[39],c56[40],s56[39]);


full_add fa56_40(s55[41],c55[41],andpr58[40],c56[41],s56[40]);


full_add fa56_41(s55[42],c55[42],andpr58[41],c56[42],s56[41]);


full_add fa56_42(s55[43],c55[43],andpr58[42],c56[43],s56[42]);


full_add fa56_43(s55[44],c55[44],andpr58[43],c56[44],s56[43]);


full_add fa56_44(s55[45],c55[45],andpr58[44],c56[45],s56[44]);


full_add fa56_45(s55[46],c55[46],andpr58[45],c56[46],s56[45]);


full_add fa56_46(s55[47],c55[47],andpr58[46],c56[47],s56[46]);


full_add fa56_47(s55[48],c55[48],andpr58[47],c56[48],s56[47]);


full_add fa56_48(s55[49],c55[49],andpr58[48],c56[49],s56[48]);


full_add fa56_49(s55[50],c55[50],andpr58[49],c56[50],s56[49]);


full_add fa56_50(s55[51],c55[51],andpr58[50],c56[51],s56[50]);


full_add fa56_51(s55[52],c55[52],andpr58[51],c56[52],s56[51]);


full_add fa56_52(s55[53],c55[53],andpr58[52],c56[53],s56[52]);


full_add fa56_53(s55[54],c55[54],andpr58[53],c56[54],s56[53]);


full_add fa56_54(s55[55],c55[55],andpr58[54],c56[55],s56[54]);


full_add fa56_55(s55[56],c55[56],andpr58[55],c56[56],s56[55]);


full_add fa56_56(s55[57],c55[57],andpr58[56],c56[57],s56[56]);


full_add fa56_57(s55[58],c55[58],andpr58[57],c56[58],s56[57]);


full_add fa56_58(s55[59],c55[59],andpr58[58],c56[59],s56[58]);


full_add fa56_59(s55[60],c55[60],andpr58[59],c56[60],s56[59]);


full_add fa56_60(s55[61],c55[61],andpr58[60],c56[61],s56[60]);


full_add fa56_61(s55[62],c55[62],andpr58[61],c56[62],s56[61]);


full_add fa56_62(si[56],c55[63],andpr58[62],c56[63],s56[62]);



half_adder ha57(s56[0],c56[0],c57[0],p[57]);


full_add fa57_0(s56[1],c56[1],andpr59[0],c57[1],s57[0]);


full_add fa57_1(s56[2],c56[2],andpr59[1],c57[2],s57[1]);


full_add fa57_2(s56[3],c56[3],andpr59[2],c57[3],s57[2]);


full_add fa57_3(s56[4],c56[4],andpr59[3],c57[4],s57[3]);


full_add fa57_4(s56[5],c56[5],andpr59[4],c57[5],s57[4]);


full_add fa57_5(s56[6],c56[6],andpr59[5],c57[6],s57[5]);


full_add fa57_6(s56[7],c56[7],andpr59[6],c57[7],s57[6]);


full_add fa57_7(s56[8],c56[8],andpr59[7],c57[8],s57[7]);


full_add fa57_8(s56[9],c56[9],andpr59[8],c57[9],s57[8]);


full_add fa57_9(s56[10],c56[10],andpr59[9],c57[10],s57[9]);


full_add fa57_10(s56[11],c56[11],andpr59[10],c57[11],s57[10]);


full_add fa57_11(s56[12],c56[12],andpr59[11],c57[12],s57[11]);


full_add fa57_12(s56[13],c56[13],andpr59[12],c57[13],s57[12]);


full_add fa57_13(s56[14],c56[14],andpr59[13],c57[14],s57[13]);


full_add fa57_14(s56[15],c56[15],andpr59[14],c57[15],s57[14]);


full_add fa57_15(s56[16],c56[16],andpr59[15],c57[16],s57[15]);


full_add fa57_16(s56[17],c56[17],andpr59[16],c57[17],s57[16]);


full_add fa57_17(s56[18],c56[18],andpr59[17],c57[18],s57[17]);


full_add fa57_18(s56[19],c56[19],andpr59[18],c57[19],s57[18]);


full_add fa57_19(s56[20],c56[20],andpr59[19],c57[20],s57[19]);


full_add fa57_20(s56[21],c56[21],andpr59[20],c57[21],s57[20]);


full_add fa57_21(s56[22],c56[22],andpr59[21],c57[22],s57[21]);


full_add fa57_22(s56[23],c56[23],andpr59[22],c57[23],s57[22]);


full_add fa57_23(s56[24],c56[24],andpr59[23],c57[24],s57[23]);


full_add fa57_24(s56[25],c56[25],andpr59[24],c57[25],s57[24]);


full_add fa57_25(s56[26],c56[26],andpr59[25],c57[26],s57[25]);


full_add fa57_26(s56[27],c56[27],andpr59[26],c57[27],s57[26]);


full_add fa57_27(s56[28],c56[28],andpr59[27],c57[28],s57[27]);


full_add fa57_28(s56[29],c56[29],andpr59[28],c57[29],s57[28]);


full_add fa57_29(s56[30],c56[30],andpr59[29],c57[30],s57[29]);


full_add fa57_30(s56[31],c56[31],andpr59[30],c57[31],s57[30]);


full_add fa57_31(s56[32],c56[32],andpr59[31],c57[32],s57[31]);


full_add fa57_32(s56[33],c56[33],andpr59[32],c57[33],s57[32]);


full_add fa57_33(s56[34],c56[34],andpr59[33],c57[34],s57[33]);


full_add fa57_34(s56[35],c56[35],andpr59[34],c57[35],s57[34]);


full_add fa57_35(s56[36],c56[36],andpr59[35],c57[36],s57[35]);


full_add fa57_36(s56[37],c56[37],andpr59[36],c57[37],s57[36]);


full_add fa57_37(s56[38],c56[38],andpr59[37],c57[38],s57[37]);


full_add fa57_38(s56[39],c56[39],andpr59[38],c57[39],s57[38]);


full_add fa57_39(s56[40],c56[40],andpr59[39],c57[40],s57[39]);


full_add fa57_40(s56[41],c56[41],andpr59[40],c57[41],s57[40]);


full_add fa57_41(s56[42],c56[42],andpr59[41],c57[42],s57[41]);


full_add fa57_42(s56[43],c56[43],andpr59[42],c57[43],s57[42]);


full_add fa57_43(s56[44],c56[44],andpr59[43],c57[44],s57[43]);


full_add fa57_44(s56[45],c56[45],andpr59[44],c57[45],s57[44]);


full_add fa57_45(s56[46],c56[46],andpr59[45],c57[46],s57[45]);


full_add fa57_46(s56[47],c56[47],andpr59[46],c57[47],s57[46]);


full_add fa57_47(s56[48],c56[48],andpr59[47],c57[48],s57[47]);


full_add fa57_48(s56[49],c56[49],andpr59[48],c57[49],s57[48]);


full_add fa57_49(s56[50],c56[50],andpr59[49],c57[50],s57[49]);


full_add fa57_50(s56[51],c56[51],andpr59[50],c57[51],s57[50]);


full_add fa57_51(s56[52],c56[52],andpr59[51],c57[52],s57[51]);


full_add fa57_52(s56[53],c56[53],andpr59[52],c57[53],s57[52]);


full_add fa57_53(s56[54],c56[54],andpr59[53],c57[54],s57[53]);


full_add fa57_54(s56[55],c56[55],andpr59[54],c57[55],s57[54]);


full_add fa57_55(s56[56],c56[56],andpr59[55],c57[56],s57[55]);


full_add fa57_56(s56[57],c56[57],andpr59[56],c57[57],s57[56]);


full_add fa57_57(s56[58],c56[58],andpr59[57],c57[58],s57[57]);


full_add fa57_58(s56[59],c56[59],andpr59[58],c57[59],s57[58]);


full_add fa57_59(s56[60],c56[60],andpr59[59],c57[60],s57[59]);


full_add fa57_60(s56[61],c56[61],andpr59[60],c57[61],s57[60]);


full_add fa57_61(s56[62],c56[62],andpr59[61],c57[62],s57[61]);


full_add fa57_62(si[57],c56[63],andpr59[62],c57[63],s57[62]);



half_adder ha58(s57[0],c57[0],c58[0],p[58]);


full_add fa58_0(s57[1],c57[1],andpr60[0],c58[1],s58[0]);


full_add fa58_1(s57[2],c57[2],andpr60[1],c58[2],s58[1]);


full_add fa58_2(s57[3],c57[3],andpr60[2],c58[3],s58[2]);


full_add fa58_3(s57[4],c57[4],andpr60[3],c58[4],s58[3]);


full_add fa58_4(s57[5],c57[5],andpr60[4],c58[5],s58[4]);


full_add fa58_5(s57[6],c57[6],andpr60[5],c58[6],s58[5]);


full_add fa58_6(s57[7],c57[7],andpr60[6],c58[7],s58[6]);


full_add fa58_7(s57[8],c57[8],andpr60[7],c58[8],s58[7]);


full_add fa58_8(s57[9],c57[9],andpr60[8],c58[9],s58[8]);


full_add fa58_9(s57[10],c57[10],andpr60[9],c58[10],s58[9]);


full_add fa58_10(s57[11],c57[11],andpr60[10],c58[11],s58[10]);


full_add fa58_11(s57[12],c57[12],andpr60[11],c58[12],s58[11]);


full_add fa58_12(s57[13],c57[13],andpr60[12],c58[13],s58[12]);


full_add fa58_13(s57[14],c57[14],andpr60[13],c58[14],s58[13]);


full_add fa58_14(s57[15],c57[15],andpr60[14],c58[15],s58[14]);


full_add fa58_15(s57[16],c57[16],andpr60[15],c58[16],s58[15]);


full_add fa58_16(s57[17],c57[17],andpr60[16],c58[17],s58[16]);


full_add fa58_17(s57[18],c57[18],andpr60[17],c58[18],s58[17]);


full_add fa58_18(s57[19],c57[19],andpr60[18],c58[19],s58[18]);


full_add fa58_19(s57[20],c57[20],andpr60[19],c58[20],s58[19]);


full_add fa58_20(s57[21],c57[21],andpr60[20],c58[21],s58[20]);


full_add fa58_21(s57[22],c57[22],andpr60[21],c58[22],s58[21]);


full_add fa58_22(s57[23],c57[23],andpr60[22],c58[23],s58[22]);


full_add fa58_23(s57[24],c57[24],andpr60[23],c58[24],s58[23]);


full_add fa58_24(s57[25],c57[25],andpr60[24],c58[25],s58[24]);


full_add fa58_25(s57[26],c57[26],andpr60[25],c58[26],s58[25]);


full_add fa58_26(s57[27],c57[27],andpr60[26],c58[27],s58[26]);


full_add fa58_27(s57[28],c57[28],andpr60[27],c58[28],s58[27]);


full_add fa58_28(s57[29],c57[29],andpr60[28],c58[29],s58[28]);


full_add fa58_29(s57[30],c57[30],andpr60[29],c58[30],s58[29]);


full_add fa58_30(s57[31],c57[31],andpr60[30],c58[31],s58[30]);


full_add fa58_31(s57[32],c57[32],andpr60[31],c58[32],s58[31]);


full_add fa58_32(s57[33],c57[33],andpr60[32],c58[33],s58[32]);


full_add fa58_33(s57[34],c57[34],andpr60[33],c58[34],s58[33]);


full_add fa58_34(s57[35],c57[35],andpr60[34],c58[35],s58[34]);


full_add fa58_35(s57[36],c57[36],andpr60[35],c58[36],s58[35]);


full_add fa58_36(s57[37],c57[37],andpr60[36],c58[37],s58[36]);


full_add fa58_37(s57[38],c57[38],andpr60[37],c58[38],s58[37]);


full_add fa58_38(s57[39],c57[39],andpr60[38],c58[39],s58[38]);


full_add fa58_39(s57[40],c57[40],andpr60[39],c58[40],s58[39]);


full_add fa58_40(s57[41],c57[41],andpr60[40],c58[41],s58[40]);


full_add fa58_41(s57[42],c57[42],andpr60[41],c58[42],s58[41]);


full_add fa58_42(s57[43],c57[43],andpr60[42],c58[43],s58[42]);


full_add fa58_43(s57[44],c57[44],andpr60[43],c58[44],s58[43]);


full_add fa58_44(s57[45],c57[45],andpr60[44],c58[45],s58[44]);


full_add fa58_45(s57[46],c57[46],andpr60[45],c58[46],s58[45]);


full_add fa58_46(s57[47],c57[47],andpr60[46],c58[47],s58[46]);


full_add fa58_47(s57[48],c57[48],andpr60[47],c58[48],s58[47]);


full_add fa58_48(s57[49],c57[49],andpr60[48],c58[49],s58[48]);


full_add fa58_49(s57[50],c57[50],andpr60[49],c58[50],s58[49]);


full_add fa58_50(s57[51],c57[51],andpr60[50],c58[51],s58[50]);


full_add fa58_51(s57[52],c57[52],andpr60[51],c58[52],s58[51]);


full_add fa58_52(s57[53],c57[53],andpr60[52],c58[53],s58[52]);


full_add fa58_53(s57[54],c57[54],andpr60[53],c58[54],s58[53]);


full_add fa58_54(s57[55],c57[55],andpr60[54],c58[55],s58[54]);


full_add fa58_55(s57[56],c57[56],andpr60[55],c58[56],s58[55]);


full_add fa58_56(s57[57],c57[57],andpr60[56],c58[57],s58[56]);


full_add fa58_57(s57[58],c57[58],andpr60[57],c58[58],s58[57]);


full_add fa58_58(s57[59],c57[59],andpr60[58],c58[59],s58[58]);


full_add fa58_59(s57[60],c57[60],andpr60[59],c58[60],s58[59]);


full_add fa58_60(s57[61],c57[61],andpr60[60],c58[61],s58[60]);


full_add fa58_61(s57[62],c57[62],andpr60[61],c58[62],s58[61]);


full_add fa58_62(si[58],c57[63],andpr60[62],c58[63],s58[62]);



half_adder ha59(s58[0],c58[0],c59[0],p[59]);


full_add fa59_0(s58[1],c58[1],andpr61[0],c59[1],s59[0]);


full_add fa59_1(s58[2],c58[2],andpr61[1],c59[2],s59[1]);


full_add fa59_2(s58[3],c58[3],andpr61[2],c59[3],s59[2]);


full_add fa59_3(s58[4],c58[4],andpr61[3],c59[4],s59[3]);


full_add fa59_4(s58[5],c58[5],andpr61[4],c59[5],s59[4]);


full_add fa59_5(s58[6],c58[6],andpr61[5],c59[6],s59[5]);


full_add fa59_6(s58[7],c58[7],andpr61[6],c59[7],s59[6]);


full_add fa59_7(s58[8],c58[8],andpr61[7],c59[8],s59[7]);


full_add fa59_8(s58[9],c58[9],andpr61[8],c59[9],s59[8]);


full_add fa59_9(s58[10],c58[10],andpr61[9],c59[10],s59[9]);


full_add fa59_10(s58[11],c58[11],andpr61[10],c59[11],s59[10]);


full_add fa59_11(s58[12],c58[12],andpr61[11],c59[12],s59[11]);


full_add fa59_12(s58[13],c58[13],andpr61[12],c59[13],s59[12]);


full_add fa59_13(s58[14],c58[14],andpr61[13],c59[14],s59[13]);


full_add fa59_14(s58[15],c58[15],andpr61[14],c59[15],s59[14]);


full_add fa59_15(s58[16],c58[16],andpr61[15],c59[16],s59[15]);


full_add fa59_16(s58[17],c58[17],andpr61[16],c59[17],s59[16]);


full_add fa59_17(s58[18],c58[18],andpr61[17],c59[18],s59[17]);


full_add fa59_18(s58[19],c58[19],andpr61[18],c59[19],s59[18]);


full_add fa59_19(s58[20],c58[20],andpr61[19],c59[20],s59[19]);


full_add fa59_20(s58[21],c58[21],andpr61[20],c59[21],s59[20]);


full_add fa59_21(s58[22],c58[22],andpr61[21],c59[22],s59[21]);


full_add fa59_22(s58[23],c58[23],andpr61[22],c59[23],s59[22]);


full_add fa59_23(s58[24],c58[24],andpr61[23],c59[24],s59[23]);


full_add fa59_24(s58[25],c58[25],andpr61[24],c59[25],s59[24]);


full_add fa59_25(s58[26],c58[26],andpr61[25],c59[26],s59[25]);


full_add fa59_26(s58[27],c58[27],andpr61[26],c59[27],s59[26]);


full_add fa59_27(s58[28],c58[28],andpr61[27],c59[28],s59[27]);


full_add fa59_28(s58[29],c58[29],andpr61[28],c59[29],s59[28]);


full_add fa59_29(s58[30],c58[30],andpr61[29],c59[30],s59[29]);


full_add fa59_30(s58[31],c58[31],andpr61[30],c59[31],s59[30]);


full_add fa59_31(s58[32],c58[32],andpr61[31],c59[32],s59[31]);


full_add fa59_32(s58[33],c58[33],andpr61[32],c59[33],s59[32]);


full_add fa59_33(s58[34],c58[34],andpr61[33],c59[34],s59[33]);


full_add fa59_34(s58[35],c58[35],andpr61[34],c59[35],s59[34]);


full_add fa59_35(s58[36],c58[36],andpr61[35],c59[36],s59[35]);


full_add fa59_36(s58[37],c58[37],andpr61[36],c59[37],s59[36]);


full_add fa59_37(s58[38],c58[38],andpr61[37],c59[38],s59[37]);


full_add fa59_38(s58[39],c58[39],andpr61[38],c59[39],s59[38]);


full_add fa59_39(s58[40],c58[40],andpr61[39],c59[40],s59[39]);


full_add fa59_40(s58[41],c58[41],andpr61[40],c59[41],s59[40]);


full_add fa59_41(s58[42],c58[42],andpr61[41],c59[42],s59[41]);


full_add fa59_42(s58[43],c58[43],andpr61[42],c59[43],s59[42]);


full_add fa59_43(s58[44],c58[44],andpr61[43],c59[44],s59[43]);


full_add fa59_44(s58[45],c58[45],andpr61[44],c59[45],s59[44]);


full_add fa59_45(s58[46],c58[46],andpr61[45],c59[46],s59[45]);


full_add fa59_46(s58[47],c58[47],andpr61[46],c59[47],s59[46]);


full_add fa59_47(s58[48],c58[48],andpr61[47],c59[48],s59[47]);


full_add fa59_48(s58[49],c58[49],andpr61[48],c59[49],s59[48]);


full_add fa59_49(s58[50],c58[50],andpr61[49],c59[50],s59[49]);


full_add fa59_50(s58[51],c58[51],andpr61[50],c59[51],s59[50]);


full_add fa59_51(s58[52],c58[52],andpr61[51],c59[52],s59[51]);


full_add fa59_52(s58[53],c58[53],andpr61[52],c59[53],s59[52]);


full_add fa59_53(s58[54],c58[54],andpr61[53],c59[54],s59[53]);


full_add fa59_54(s58[55],c58[55],andpr61[54],c59[55],s59[54]);


full_add fa59_55(s58[56],c58[56],andpr61[55],c59[56],s59[55]);


full_add fa59_56(s58[57],c58[57],andpr61[56],c59[57],s59[56]);


full_add fa59_57(s58[58],c58[58],andpr61[57],c59[58],s59[57]);


full_add fa59_58(s58[59],c58[59],andpr61[58],c59[59],s59[58]);


full_add fa59_59(s58[60],c58[60],andpr61[59],c59[60],s59[59]);


full_add fa59_60(s58[61],c58[61],andpr61[60],c59[61],s59[60]);


full_add fa59_61(s58[62],c58[62],andpr61[61],c59[62],s59[61]);


full_add fa59_62(si[59],c58[63],andpr61[62],c59[63],s59[62]);



half_adder ha60(s59[0],c59[0],c60[0],p[60]);


full_add fa60_0(s59[1],c59[1],andpr62[0],c60[1],s60[0]);


full_add fa60_1(s59[2],c59[2],andpr62[1],c60[2],s60[1]);


full_add fa60_2(s59[3],c59[3],andpr62[2],c60[3],s60[2]);


full_add fa60_3(s59[4],c59[4],andpr62[3],c60[4],s60[3]);


full_add fa60_4(s59[5],c59[5],andpr62[4],c60[5],s60[4]);


full_add fa60_5(s59[6],c59[6],andpr62[5],c60[6],s60[5]);


full_add fa60_6(s59[7],c59[7],andpr62[6],c60[7],s60[6]);


full_add fa60_7(s59[8],c59[8],andpr62[7],c60[8],s60[7]);


full_add fa60_8(s59[9],c59[9],andpr62[8],c60[9],s60[8]);


full_add fa60_9(s59[10],c59[10],andpr62[9],c60[10],s60[9]);


full_add fa60_10(s59[11],c59[11],andpr62[10],c60[11],s60[10]);


full_add fa60_11(s59[12],c59[12],andpr62[11],c60[12],s60[11]);


full_add fa60_12(s59[13],c59[13],andpr62[12],c60[13],s60[12]);


full_add fa60_13(s59[14],c59[14],andpr62[13],c60[14],s60[13]);


full_add fa60_14(s59[15],c59[15],andpr62[14],c60[15],s60[14]);


full_add fa60_15(s59[16],c59[16],andpr62[15],c60[16],s60[15]);


full_add fa60_16(s59[17],c59[17],andpr62[16],c60[17],s60[16]);


full_add fa60_17(s59[18],c59[18],andpr62[17],c60[18],s60[17]);


full_add fa60_18(s59[19],c59[19],andpr62[18],c60[19],s60[18]);


full_add fa60_19(s59[20],c59[20],andpr62[19],c60[20],s60[19]);


full_add fa60_20(s59[21],c59[21],andpr62[20],c60[21],s60[20]);


full_add fa60_21(s59[22],c59[22],andpr62[21],c60[22],s60[21]);


full_add fa60_22(s59[23],c59[23],andpr62[22],c60[23],s60[22]);


full_add fa60_23(s59[24],c59[24],andpr62[23],c60[24],s60[23]);


full_add fa60_24(s59[25],c59[25],andpr62[24],c60[25],s60[24]);


full_add fa60_25(s59[26],c59[26],andpr62[25],c60[26],s60[25]);


full_add fa60_26(s59[27],c59[27],andpr62[26],c60[27],s60[26]);


full_add fa60_27(s59[28],c59[28],andpr62[27],c60[28],s60[27]);


full_add fa60_28(s59[29],c59[29],andpr62[28],c60[29],s60[28]);


full_add fa60_29(s59[30],c59[30],andpr62[29],c60[30],s60[29]);


full_add fa60_30(s59[31],c59[31],andpr62[30],c60[31],s60[30]);


full_add fa60_31(s59[32],c59[32],andpr62[31],c60[32],s60[31]);


full_add fa60_32(s59[33],c59[33],andpr62[32],c60[33],s60[32]);


full_add fa60_33(s59[34],c59[34],andpr62[33],c60[34],s60[33]);


full_add fa60_34(s59[35],c59[35],andpr62[34],c60[35],s60[34]);


full_add fa60_35(s59[36],c59[36],andpr62[35],c60[36],s60[35]);


full_add fa60_36(s59[37],c59[37],andpr62[36],c60[37],s60[36]);


full_add fa60_37(s59[38],c59[38],andpr62[37],c60[38],s60[37]);


full_add fa60_38(s59[39],c59[39],andpr62[38],c60[39],s60[38]);


full_add fa60_39(s59[40],c59[40],andpr62[39],c60[40],s60[39]);


full_add fa60_40(s59[41],c59[41],andpr62[40],c60[41],s60[40]);


full_add fa60_41(s59[42],c59[42],andpr62[41],c60[42],s60[41]);


full_add fa60_42(s59[43],c59[43],andpr62[42],c60[43],s60[42]);


full_add fa60_43(s59[44],c59[44],andpr62[43],c60[44],s60[43]);


full_add fa60_44(s59[45],c59[45],andpr62[44],c60[45],s60[44]);


full_add fa60_45(s59[46],c59[46],andpr62[45],c60[46],s60[45]);


full_add fa60_46(s59[47],c59[47],andpr62[46],c60[47],s60[46]);


full_add fa60_47(s59[48],c59[48],andpr62[47],c60[48],s60[47]);


full_add fa60_48(s59[49],c59[49],andpr62[48],c60[49],s60[48]);


full_add fa60_49(s59[50],c59[50],andpr62[49],c60[50],s60[49]);


full_add fa60_50(s59[51],c59[51],andpr62[50],c60[51],s60[50]);


full_add fa60_51(s59[52],c59[52],andpr62[51],c60[52],s60[51]);


full_add fa60_52(s59[53],c59[53],andpr62[52],c60[53],s60[52]);


full_add fa60_53(s59[54],c59[54],andpr62[53],c60[54],s60[53]);


full_add fa60_54(s59[55],c59[55],andpr62[54],c60[55],s60[54]);


full_add fa60_55(s59[56],c59[56],andpr62[55],c60[56],s60[55]);


full_add fa60_56(s59[57],c59[57],andpr62[56],c60[57],s60[56]);


full_add fa60_57(s59[58],c59[58],andpr62[57],c60[58],s60[57]);


full_add fa60_58(s59[59],c59[59],andpr62[58],c60[59],s60[58]);


full_add fa60_59(s59[60],c59[60],andpr62[59],c60[60],s60[59]);


full_add fa60_60(s59[61],c59[61],andpr62[60],c60[61],s60[60]);


full_add fa60_61(s59[62],c59[62],andpr62[61],c60[62],s60[61]);


full_add fa60_62(si[60],c59[63],andpr62[62],c60[63],s60[62]);



half_adder ha61(s60[0],c60[0],c61[0],p[61]);


full_add fa61_0(s60[1],c60[1],andpr63[0],c61[1],s61[0]);


full_add fa61_1(s60[2],c60[2],andpr63[1],c61[2],s61[1]);


full_add fa61_2(s60[3],c60[3],andpr63[2],c61[3],s61[2]);


full_add fa61_3(s60[4],c60[4],andpr63[3],c61[4],s61[3]);


full_add fa61_4(s60[5],c60[5],andpr63[4],c61[5],s61[4]);


full_add fa61_5(s60[6],c60[6],andpr63[5],c61[6],s61[5]);


full_add fa61_6(s60[7],c60[7],andpr63[6],c61[7],s61[6]);


full_add fa61_7(s60[8],c60[8],andpr63[7],c61[8],s61[7]);


full_add fa61_8(s60[9],c60[9],andpr63[8],c61[9],s61[8]);


full_add fa61_9(s60[10],c60[10],andpr63[9],c61[10],s61[9]);


full_add fa61_10(s60[11],c60[11],andpr63[10],c61[11],s61[10]);


full_add fa61_11(s60[12],c60[12],andpr63[11],c61[12],s61[11]);


full_add fa61_12(s60[13],c60[13],andpr63[12],c61[13],s61[12]);


full_add fa61_13(s60[14],c60[14],andpr63[13],c61[14],s61[13]);


full_add fa61_14(s60[15],c60[15],andpr63[14],c61[15],s61[14]);


full_add fa61_15(s60[16],c60[16],andpr63[15],c61[16],s61[15]);


full_add fa61_16(s60[17],c60[17],andpr63[16],c61[17],s61[16]);


full_add fa61_17(s60[18],c60[18],andpr63[17],c61[18],s61[17]);


full_add fa61_18(s60[19],c60[19],andpr63[18],c61[19],s61[18]);


full_add fa61_19(s60[20],c60[20],andpr63[19],c61[20],s61[19]);


full_add fa61_20(s60[21],c60[21],andpr63[20],c61[21],s61[20]);


full_add fa61_21(s60[22],c60[22],andpr63[21],c61[22],s61[21]);


full_add fa61_22(s60[23],c60[23],andpr63[22],c61[23],s61[22]);


full_add fa61_23(s60[24],c60[24],andpr63[23],c61[24],s61[23]);


full_add fa61_24(s60[25],c60[25],andpr63[24],c61[25],s61[24]);


full_add fa61_25(s60[26],c60[26],andpr63[25],c61[26],s61[25]);


full_add fa61_26(s60[27],c60[27],andpr63[26],c61[27],s61[26]);


full_add fa61_27(s60[28],c60[28],andpr63[27],c61[28],s61[27]);


full_add fa61_28(s60[29],c60[29],andpr63[28],c61[29],s61[28]);


full_add fa61_29(s60[30],c60[30],andpr63[29],c61[30],s61[29]);


full_add fa61_30(s60[31],c60[31],andpr63[30],c61[31],s61[30]);


full_add fa61_31(s60[32],c60[32],andpr63[31],c61[32],s61[31]);


full_add fa61_32(s60[33],c60[33],andpr63[32],c61[33],s61[32]);


full_add fa61_33(s60[34],c60[34],andpr63[33],c61[34],s61[33]);


full_add fa61_34(s60[35],c60[35],andpr63[34],c61[35],s61[34]);


full_add fa61_35(s60[36],c60[36],andpr63[35],c61[36],s61[35]);


full_add fa61_36(s60[37],c60[37],andpr63[36],c61[37],s61[36]);


full_add fa61_37(s60[38],c60[38],andpr63[37],c61[38],s61[37]);


full_add fa61_38(s60[39],c60[39],andpr63[38],c61[39],s61[38]);


full_add fa61_39(s60[40],c60[40],andpr63[39],c61[40],s61[39]);


full_add fa61_40(s60[41],c60[41],andpr63[40],c61[41],s61[40]);


full_add fa61_41(s60[42],c60[42],andpr63[41],c61[42],s61[41]);


full_add fa61_42(s60[43],c60[43],andpr63[42],c61[43],s61[42]);


full_add fa61_43(s60[44],c60[44],andpr63[43],c61[44],s61[43]);


full_add fa61_44(s60[45],c60[45],andpr63[44],c61[45],s61[44]);


full_add fa61_45(s60[46],c60[46],andpr63[45],c61[46],s61[45]);


full_add fa61_46(s60[47],c60[47],andpr63[46],c61[47],s61[46]);


full_add fa61_47(s60[48],c60[48],andpr63[47],c61[48],s61[47]);


full_add fa61_48(s60[49],c60[49],andpr63[48],c61[49],s61[48]);


full_add fa61_49(s60[50],c60[50],andpr63[49],c61[50],s61[49]);


full_add fa61_50(s60[51],c60[51],andpr63[50],c61[51],s61[50]);


full_add fa61_51(s60[52],c60[52],andpr63[51],c61[52],s61[51]);


full_add fa61_52(s60[53],c60[53],andpr63[52],c61[53],s61[52]);


full_add fa61_53(s60[54],c60[54],andpr63[53],c61[54],s61[53]);


full_add fa61_54(s60[55],c60[55],andpr63[54],c61[55],s61[54]);


full_add fa61_55(s60[56],c60[56],andpr63[55],c61[56],s61[55]);


full_add fa61_56(s60[57],c60[57],andpr63[56],c61[57],s61[56]);


full_add fa61_57(s60[58],c60[58],andpr63[57],c61[58],s61[57]);


full_add fa61_58(s60[59],c60[59],andpr63[58],c61[59],s61[58]);


full_add fa61_59(s60[60],c60[60],andpr63[59],c61[60],s61[59]);


full_add fa61_60(s60[61],c60[61],andpr63[60],c61[61],s61[60]);


full_add fa61_61(s60[62],c60[62],andpr63[61],c61[62],s61[61]);


full_add fa61_62(si[61],c60[63],andpr63[62],c61[63],s61[62]);



half_adder ha62(s61[0],c61[0],c62[0],p[62]);


full_add fa62_0(s61[1],c61[1],andpr64[0],c62[1],s62[0]);


full_add fa62_1(s61[2],c61[2],andpr64[1],c62[2],s62[1]);


full_add fa62_2(s61[3],c61[3],andpr64[2],c62[3],s62[2]);


full_add fa62_3(s61[4],c61[4],andpr64[3],c62[4],s62[3]);


full_add fa62_4(s61[5],c61[5],andpr64[4],c62[5],s62[4]);


full_add fa62_5(s61[6],c61[6],andpr64[5],c62[6],s62[5]);


full_add fa62_6(s61[7],c61[7],andpr64[6],c62[7],s62[6]);


full_add fa62_7(s61[8],c61[8],andpr64[7],c62[8],s62[7]);


full_add fa62_8(s61[9],c61[9],andpr64[8],c62[9],s62[8]);


full_add fa62_9(s61[10],c61[10],andpr64[9],c62[10],s62[9]);


full_add fa62_10(s61[11],c61[11],andpr64[10],c62[11],s62[10]);


full_add fa62_11(s61[12],c61[12],andpr64[11],c62[12],s62[11]);


full_add fa62_12(s61[13],c61[13],andpr64[12],c62[13],s62[12]);


full_add fa62_13(s61[14],c61[14],andpr64[13],c62[14],s62[13]);


full_add fa62_14(s61[15],c61[15],andpr64[14],c62[15],s62[14]);


full_add fa62_15(s61[16],c61[16],andpr64[15],c62[16],s62[15]);


full_add fa62_16(s61[17],c61[17],andpr64[16],c62[17],s62[16]);


full_add fa62_17(s61[18],c61[18],andpr64[17],c62[18],s62[17]);


full_add fa62_18(s61[19],c61[19],andpr64[18],c62[19],s62[18]);


full_add fa62_19(s61[20],c61[20],andpr64[19],c62[20],s62[19]);


full_add fa62_20(s61[21],c61[21],andpr64[20],c62[21],s62[20]);


full_add fa62_21(s61[22],c61[22],andpr64[21],c62[22],s62[21]);


full_add fa62_22(s61[23],c61[23],andpr64[22],c62[23],s62[22]);


full_add fa62_23(s61[24],c61[24],andpr64[23],c62[24],s62[23]);


full_add fa62_24(s61[25],c61[25],andpr64[24],c62[25],s62[24]);


full_add fa62_25(s61[26],c61[26],andpr64[25],c62[26],s62[25]);


full_add fa62_26(s61[27],c61[27],andpr64[26],c62[27],s62[26]);


full_add fa62_27(s61[28],c61[28],andpr64[27],c62[28],s62[27]);


full_add fa62_28(s61[29],c61[29],andpr64[28],c62[29],s62[28]);


full_add fa62_29(s61[30],c61[30],andpr64[29],c62[30],s62[29]);


full_add fa62_30(s61[31],c61[31],andpr64[30],c62[31],s62[30]);


full_add fa62_31(s61[32],c61[32],andpr64[31],c62[32],s62[31]);


full_add fa62_32(s61[33],c61[33],andpr64[32],c62[33],s62[32]);


full_add fa62_33(s61[34],c61[34],andpr64[33],c62[34],s62[33]);


full_add fa62_34(s61[35],c61[35],andpr64[34],c62[35],s62[34]);


full_add fa62_35(s61[36],c61[36],andpr64[35],c62[36],s62[35]);


full_add fa62_36(s61[37],c61[37],andpr64[36],c62[37],s62[36]);


full_add fa62_37(s61[38],c61[38],andpr64[37],c62[38],s62[37]);


full_add fa62_38(s61[39],c61[39],andpr64[38],c62[39],s62[38]);


full_add fa62_39(s61[40],c61[40],andpr64[39],c62[40],s62[39]);


full_add fa62_40(s61[41],c61[41],andpr64[40],c62[41],s62[40]);


full_add fa62_41(s61[42],c61[42],andpr64[41],c62[42],s62[41]);


full_add fa62_42(s61[43],c61[43],andpr64[42],c62[43],s62[42]);


full_add fa62_43(s61[44],c61[44],andpr64[43],c62[44],s62[43]);


full_add fa62_44(s61[45],c61[45],andpr64[44],c62[45],s62[44]);


full_add fa62_45(s61[46],c61[46],andpr64[45],c62[46],s62[45]);


full_add fa62_46(s61[47],c61[47],andpr64[46],c62[47],s62[46]);


full_add fa62_47(s61[48],c61[48],andpr64[47],c62[48],s62[47]);


full_add fa62_48(s61[49],c61[49],andpr64[48],c62[49],s62[48]);


full_add fa62_49(s61[50],c61[50],andpr64[49],c62[50],s62[49]);


full_add fa62_50(s61[51],c61[51],andpr64[50],c62[51],s62[50]);


full_add fa62_51(s61[52],c61[52],andpr64[51],c62[52],s62[51]);


full_add fa62_52(s61[53],c61[53],andpr64[52],c62[53],s62[52]);


full_add fa62_53(s61[54],c61[54],andpr64[53],c62[54],s62[53]);


full_add fa62_54(s61[55],c61[55],andpr64[54],c62[55],s62[54]);


full_add fa62_55(s61[56],c61[56],andpr64[55],c62[56],s62[55]);


full_add fa62_56(s61[57],c61[57],andpr64[56],c62[57],s62[56]);


full_add fa62_57(s61[58],c61[58],andpr64[57],c62[58],s62[57]);


full_add fa62_58(s61[59],c61[59],andpr64[58],c62[59],s62[58]);


full_add fa62_59(s61[60],c61[60],andpr64[59],c62[60],s62[59]);


full_add fa62_60(s61[61],c61[61],andpr64[60],c62[61],s62[60]);


full_add fa62_61(s61[62],c61[62],andpr64[61],c62[62],s62[61]);


full_add fa62_62(si[62],c61[63],andpr64[62],c62[63],s62[62]);



//last layer
full_add fad63_62(s62[0],c62[0],b[63],c63[0],p[63]);


full_add fad63_63(s62[1],c62[1],c63[0],c63[1],p[64]);


full_add fad63_64(s62[2],c62[2],c63[1],c63[2],p[65]);


full_add fad63_65(s62[3],c62[3],c63[2],c63[3],p[66]);


full_add fad63_66(s62[4],c62[4],c63[3],c63[4],p[67]);


full_add fad63_67(s62[5],c62[5],c63[4],c63[5],p[68]);


full_add fad63_68(s62[6],c62[6],c63[5],c63[6],p[69]);


full_add fad63_69(s62[7],c62[7],c63[6],c63[7],p[70]);


full_add fad63_70(s62[8],c62[8],c63[7],c63[8],p[71]);


full_add fad63_71(s62[9],c62[9],c63[8],c63[9],p[72]);


full_add fad63_72(s62[10],c62[10],c63[9],c63[10],p[73]);


full_add fad63_73(s62[11],c62[11],c63[10],c63[11],p[74]);


full_add fad63_74(s62[12],c62[12],c63[11],c63[12],p[75]);


full_add fad63_75(s62[13],c62[13],c63[12],c63[13],p[76]);


full_add fad63_76(s62[14],c62[14],c63[13],c63[14],p[77]);


full_add fad63_77(s62[15],c62[15],c63[14],c63[15],p[78]);


full_add fad63_78(s62[16],c62[16],c63[15],c63[16],p[79]);


full_add fad63_79(s62[17],c62[17],c63[16],c63[17],p[80]);


full_add fad63_80(s62[18],c62[18],c63[17],c63[18],p[81]);


full_add fad63_81(s62[19],c62[19],c63[18],c63[19],p[82]);


full_add fad63_82(s62[20],c62[20],c63[19],c63[20],p[83]);


full_add fad63_83(s62[21],c62[21],c63[20],c63[21],p[84]);


full_add fad63_84(s62[22],c62[22],c63[21],c63[22],p[85]);


full_add fad63_85(s62[23],c62[23],c63[22],c63[23],p[86]);


full_add fad63_86(s62[24],c62[24],c63[23],c63[24],p[87]);


full_add fad63_87(s62[25],c62[25],c63[24],c63[25],p[88]);


full_add fad63_88(s62[26],c62[26],c63[25],c63[26],p[89]);


full_add fad63_89(s62[27],c62[27],c63[26],c63[27],p[90]);


full_add fad63_90(s62[28],c62[28],c63[27],c63[28],p[91]);


full_add fad63_91(s62[29],c62[29],c63[28],c63[29],p[92]);


full_add fad63_92(s62[30],c62[30],c63[29],c63[30],p[93]);


full_add fad63_93(s62[31],c62[31],c63[30],c63[31],p[94]);


full_add fad63_94(s62[32],c62[32],c63[31],c63[32],p[95]);


full_add fad63_95(s62[33],c62[33],c63[32],c63[33],p[96]);


full_add fad63_96(s62[34],c62[34],c63[33],c63[34],p[97]);


full_add fad63_97(s62[35],c62[35],c63[34],c63[35],p[98]);


full_add fad63_98(s62[36],c62[36],c63[35],c63[36],p[99]);


full_add fad63_99(s62[37],c62[37],c63[36],c63[37],p[100]);


full_add fad63_100(s62[38],c62[38],c63[37],c63[38],p[101]);


full_add fad63_101(s62[39],c62[39],c63[38],c63[39],p[102]);


full_add fad63_102(s62[40],c62[40],c63[39],c63[40],p[103]);


full_add fad63_103(s62[41],c62[41],c63[40],c63[41],p[104]);


full_add fad63_104(s62[42],c62[42],c63[41],c63[42],p[105]);


full_add fad63_105(s62[43],c62[43],c63[42],c63[43],p[106]);


full_add fad63_106(s62[44],c62[44],c63[43],c63[44],p[107]);


full_add fad63_107(s62[45],c62[45],c63[44],c63[45],p[108]);


full_add fad63_108(s62[46],c62[46],c63[45],c63[46],p[109]);


full_add fad63_109(s62[47],c62[47],c63[46],c63[47],p[110]);


full_add fad63_110(s62[48],c62[48],c63[47],c63[48],p[111]);


full_add fad63_111(s62[49],c62[49],c63[48],c63[49],p[112]);


full_add fad63_112(s62[50],c62[50],c63[49],c63[50],p[113]);


full_add fad63_113(s62[51],c62[51],c63[50],c63[51],p[114]);


full_add fad63_114(s62[52],c62[52],c63[51],c63[52],p[115]);


full_add fad63_115(s62[53],c62[53],c63[52],c63[53],p[116]);


full_add fad63_116(s62[54],c62[54],c63[53],c63[54],p[117]);


full_add fad63_117(s62[55],c62[55],c63[54],c63[55],p[118]);


full_add fad63_118(s62[56],c62[56],c63[55],c63[56],p[119]);


full_add fad63_119(s62[57],c62[57],c63[56],c63[57],p[120]);


full_add fad63_120(s62[58],c62[58],c63[57],c63[58],p[121]);


full_add fad63_121(s62[59],c62[59],c63[58],c63[59],p[122]);


full_add fad63_122(s62[60],c62[60],c63[59],c63[60],p[123]);


full_add fad63_123(s62[61],c62[61],c63[60],c63[61],p[124]);


full_add fad63_124(s62[62],c62[62],c63[61],c63[62],p[125]);


full_add fad63_125(si[63],c62[63],c63[62],c63[63],p[126]);
half_adder ha64(c63[63],1'b1,c,p[127]);
assign p[0]=andpr1[0];

endmodule